-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_F2 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_F2 is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"00",x"00",x"71",x"C0",x"F1",x"E0",x"87",x"2C", -- 0x0000
		x"80",x"20",x"F1",x"E0",x"79",x"C2",x"07",x"0C", -- 0x0008
		x"00",x"00",x"80",x"80",x"80",x"48",x"F1",x"E0", -- 0x0010
		x"F1",x"E0",x"87",x"0E",x"80",x"00",x"08",x"00", -- 0x0018
		x"00",x"00",x"C0",x"40",x"E0",x"60",x"A4",x"24", -- 0x0020
		x"93",x"20",x"91",x"E0",x"81",x"C2",x"08",x"0C", -- 0x0028
		x"00",x"00",x"40",x"40",x"C0",x"60",x"95",x"24", -- 0x0030
		x"91",x"20",x"F1",x"E0",x"69",x"C2",x"06",x"0C", -- 0x0038
		x"00",x"00",x"31",x"00",x"31",x"80",x"21",x"C0", -- 0x0040
		x"20",x"68",x"F1",x"E0",x"F1",x"E0",x"2D",x"0E", -- 0x0048
		x"00",x"00",x"51",x"E0",x"D1",x"E0",x"85",x"A4", -- 0x0050
		x"80",x"A0",x"F1",x"A0",x"79",x"28",x"07",x"02", -- 0x0058
		x"00",x"00",x"71",x"C0",x"F1",x"E0",x"97",x"2C", -- 0x0060
		x"91",x"20",x"F1",x"60",x"69",x"42",x"06",x"04", -- 0x0068
		x"00",x"00",x"00",x"20",x"E0",x"20",x"F1",x"20", -- 0x0070
		x"1F",x"A0",x"01",x"E0",x"00",x"68",x"00",x"06", -- 0x0078
		x"00",x"00",x"60",x"C0",x"F1",x"E0",x"97",x"2C", -- 0x0080
		x"91",x"20",x"F1",x"E0",x"69",x"C2",x"06",x"0C", -- 0x0088
		x"00",x"00",x"00",x"C0",x"91",x"E0",x"91",x"2C", -- 0x0090
		x"91",x"20",x"79",x"E0",x"35",x"C2",x"03",x"0C", -- 0x0098
		x"00",x"00",x"79",x"80",x"79",x"C0",x"20",x"42", -- 0x00A0
		x"20",x"02",x"20",x"42",x"79",x"C0",x"79",x"80", -- 0x00A8
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"19",x"02", -- 0x00B0
		x"19",x"02",x"19",x"02",x"79",x"C2",x"60",x"C0", -- 0x00B8
		x"00",x"00",x"71",x"C0",x"79",x"C2",x"08",x"02", -- 0x00C0
		x"08",x"02",x"08",x"02",x"48",x"42",x"40",x"40", -- 0x00C8
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"08",x"02", -- 0x00D0
		x"08",x"02",x"08",x"02",x"79",x"C2",x"71",x"C0", -- 0x00D8
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"19",x"02", -- 0x00E0
		x"19",x"02",x"19",x"02",x"19",x"02",x"08",x"02", -- 0x00E8
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"11",x"02", -- 0x00F0
		x"11",x"02",x"11",x"02",x"11",x"02",x"00",x"02", -- 0x00F8
		x"00",x"00",x"71",x"C0",x"79",x"C2",x"08",x"02", -- 0x0100
		x"08",x"02",x"28",x"02",x"68",x"42",x"60",x"40", -- 0x0108
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"11",x"00", -- 0x0110
		x"11",x"00",x"11",x"00",x"79",x"C2",x"79",x"C2", -- 0x0118
		x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"02", -- 0x0120
		x"79",x"C2",x"79",x"C2",x"08",x"02",x"00",x"00", -- 0x0128
		x"00",x"00",x"40",x"00",x"48",x"00",x"08",x"00", -- 0x0130
		x"08",x"02",x"79",x"C2",x"71",x"C2",x"00",x"02", -- 0x0138
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"31",x"00", -- 0x0140
		x"31",x"80",x"60",x"C0",x"48",x"42",x"08",x"02", -- 0x0148
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"08",x"00", -- 0x0150
		x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00", -- 0x0158
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"00",x"C0", -- 0x0160
		x"11",x"80",x"00",x"C0",x"79",x"C2",x"79",x"C2", -- 0x0168
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"00",x"C0", -- 0x0170
		x"11",x"80",x"31",x"00",x"79",x"C2",x"79",x"C2", -- 0x0178
		x"00",x"00",x"71",x"C0",x"79",x"C2",x"08",x"02", -- 0x0180
		x"08",x"02",x"08",x"02",x"79",x"C2",x"71",x"C0", -- 0x0188
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"11",x"02", -- 0x0190
		x"11",x"02",x"11",x"02",x"11",x"C2",x"00",x"C0", -- 0x0198
		x"00",x"00",x"71",x"C0",x"79",x"C2",x"08",x"02", -- 0x01A0
		x"08",x"02",x"40",x"02",x"79",x"C2",x"39",x"C0", -- 0x01A8
		x"00",x"00",x"79",x"C2",x"79",x"C2",x"11",x"02", -- 0x01B0
		x"31",x"02",x"71",x"02",x"59",x"C2",x"08",x"C0", -- 0x01B8
		x"00",x"00",x"40",x"C0",x"59",x"C2",x"19",x"02", -- 0x01C0
		x"19",x"02",x"19",x"02",x"79",x"42",x"60",x"40", -- 0x01C8
		x"00",x"00",x"00",x"02",x"00",x"02",x"00",x"02", -- 0x01D0
		x"79",x"C2",x"79",x"C2",x"00",x"02",x"00",x"02", -- 0x01D8
		x"00",x"00",x"71",x"C2",x"79",x"C2",x"08",x"00", -- 0x01E0
		x"08",x"00",x"08",x"00",x"79",x"C2",x"71",x"C2", -- 0x01E8
		x"00",x"00",x"00",x"00",x"31",x"C2",x"71",x"C2", -- 0x01F0
		x"08",x"00",x"08",x"00",x"71",x"C2",x"31",x"C2", -- 0x01F8
		x"00",x"00",x"71",x"C2",x"79",x"C2",x"48",x"00", -- 0x0200
		x"60",x"00",x"48",x"00",x"79",x"C2",x"71",x"C2", -- 0x0208
		x"00",x"00",x"48",x"02",x"60",x"42",x"31",x"C0", -- 0x0210
		x"11",x"80",x"31",x"C0",x"60",x"42",x"48",x"02", -- 0x0218
		x"00",x"00",x"00",x"00",x"00",x"C2",x"11",x"C2", -- 0x0220
		x"79",x"00",x"79",x"00",x"11",x"C2",x"00",x"C2", -- 0x0228
		x"00",x"00",x"08",x"02",x"48",x"02",x"68",x"02", -- 0x0230
		x"39",x"02",x"19",x"82",x"08",x"C2",x"08",x"42", -- 0x0238
		x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"00", -- 0x0240
		x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0248
		x"00",x"00",x"11",x"00",x"11",x"00",x"11",x"00", -- 0x0250
		x"11",x"00",x"11",x"00",x"11",x"00",x"11",x"00", -- 0x0258
		x"00",x"00",x"71",x"40",x"79",x"C2",x"08",x"82", -- 0x0260
		x"08",x"82",x"28",x"02",x"60",x"40",x"20",x"00", -- 0x0268
		x"00",x"00",x"00",x"C0",x"00",x"C2",x"00",x"02", -- 0x0270
		x"28",x"02",x"11",x"02",x"11",x"C2",x"00",x"C0", -- 0x0278
		x"00",x"00",x"00",x"00",x"00",x"00",x"51",x"C2", -- 0x0280
		x"51",x"C2",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0288
		x"00",x"00",x"48",x"C0",x"60",x"C0",x"31",x"00", -- 0x0290
		x"11",x"80",x"60",x"C0",x"60",x"42",x"00",x"00", -- 0x0298
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02A0
		x"71",x"C0",x"79",x"C2",x"08",x"02",x"00",x"00", -- 0x02A8
		x"00",x"00",x"08",x"02",x"79",x"C2",x"71",x"C0", -- 0x02B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x02B8
		x"00",x"00",x"40",x"80",x"68",x"40",x"19",x"C2", -- 0x02C0
		x"19",x"C2",x"68",x"40",x"40",x"80",x"00",x"00", -- 0x02C8
		x"00",x"00",x"20",x"40",x"20",x"C2",x"79",x"02", -- 0x02D0
		x"79",x"02",x"20",x"C2",x"20",x"40",x"00",x"00", -- 0x02D8
		x"00",x"00",x"10",x"C0",x"31",x"EC",x"70",x"E0", -- 0x02E0
		x"F0",x"C0",x"70",x"E0",x"30",x"E0",x"10",x"C0", -- 0x02E8
		x"00",x"00",x"20",x"40",x"71",x"C2",x"20",x"40", -- 0x02F0
		x"20",x"40",x"71",x"C2",x"20",x"40",x"00",x"00", -- 0x02F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0300
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0308
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x0310
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x0318
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x0320
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x0328
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0330
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0338
		x"00",x"00",x"00",x"00",x"08",x"00",x"60",x"00", -- 0x0340
		x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0348
		x"00",x"C0",x"00",x"C0",x"00",x"C0",x"00",x"C0", -- 0x0350
		x"00",x"C0",x"00",x"C0",x"00",x"C0",x"00",x"C0", -- 0x0358
		x"00",x"00",x"11",x"00",x"11",x"00",x"71",x"C0", -- 0x0360
		x"71",x"C0",x"11",x"00",x"11",x"00",x"00",x"00", -- 0x0368
		x"00",x"00",x"00",x"00",x"48",x"C0",x"71",x"80", -- 0x0370
		x"31",x"00",x"71",x"80",x"48",x"C0",x"00",x"00", -- 0x0378
		x"00",x"00",x"31",x"80",x"40",x"40",x"19",x"02", -- 0x0380
		x"28",x"82",x"28",x"82",x"40",x"40",x"31",x"80", -- 0x0388
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0390
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0398
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03A8
		x"00",x"00",x"11",x"E1",x"00",x"41",x"11",x"A1", -- 0x03B0
		x"00",x"00",x"71",x"00",x"08",x"00",x"71",x"00", -- 0x03B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
		x"00",x"00",x"11",x"E1",x"11",x"41",x"11",x"01", -- 0x03D0
		x"00",x"00",x"79",x"80",x"08",x"80",x"71",x"00", -- 0x03D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
		x"00",x"C0",x"0D",x"48",x"0F",x"68",x"0D",x"FC", -- 0x0400
		x"0D",x"03",x"0F",x"0E",x"0D",x"0C",x"00",x"0C", -- 0x0408
		x"68",x"30",x"5A",x"52",x"4B",x"96",x"49",x"1A", -- 0x0410
		x"48",x"12",x"68",x"34",x"4A",x"16",x"0C",x"03", -- 0x0418
		x"4C",x"00",x"6E",x"00",x"5F",x"00",x"0F",x"88", -- 0x0420
		x"01",x"4C",x"00",x"2E",x"7F",x"EE",x"0F",x"0E", -- 0x0428
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0430
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
		x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"60", -- 0x0440
		x"60",x"60",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0448
		x"00",x"00",x"10",x"00",x"10",x"00",x"00",x"00", -- 0x0450
		x"00",x"00",x"10",x"00",x"10",x"00",x"00",x"00", -- 0x0458
		x"00",x"00",x"00",x"00",x"20",x"00",x"10",x"00", -- 0x0460
		x"00",x"80",x"00",x"40",x"00",x"00",x"00",x"00", -- 0x0468
		x"00",x"00",x"10",x"00",x"10",x"00",x"10",x"00", -- 0x0470
		x"50",x"40",x"30",x"80",x"10",x"00",x"00",x"00", -- 0x0478
		x"00",x"00",x"00",x"00",x"10",x"00",x"20",x"80", -- 0x0480
		x"40",x"40",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0488
		x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"40", -- 0x0490
		x"20",x"80",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x0498
		x"00",x"00",x"00",x"00",x"20",x"80",x"20",x"80", -- 0x04A0
		x"20",x"80",x"20",x"80",x"00",x"00",x"00",x"00", -- 0x04A8
		x"00",x"00",x"20",x"40",x"10",x"80",x"70",x"E0", -- 0x04B0
		x"10",x"80",x"20",x"40",x"00",x"00",x"00",x"00", -- 0x04B8
		x"F0",x"F0",x"80",x"00",x"80",x"00",x"80",x"00", -- 0x04C0
		x"80",x"00",x"80",x"00",x"80",x"00",x"80",x"00", -- 0x04C8
		x"F0",x"F0",x"00",x"10",x"00",x"10",x"00",x"10", -- 0x04D0
		x"00",x"10",x"00",x"10",x"00",x"10",x"00",x"10", -- 0x04D8
		x"80",x"00",x"80",x"00",x"80",x"00",x"80",x"00", -- 0x04E0
		x"80",x"00",x"80",x"00",x"80",x"00",x"F0",x"F0", -- 0x04E8
		x"80",x"10",x"00",x"10",x"00",x"10",x"00",x"10", -- 0x04F0
		x"00",x"10",x"00",x"10",x"00",x"10",x"F0",x"F0", -- 0x04F8
		x"70",x"C0",x"00",x"80",x"10",x"00",x"70",x"C0", -- 0x0500
		x"00",x"00",x"70",x"00",x"50",x"00",x"70",x"00", -- 0x0508
		x"00",x"00",x"70",x"E0",x"F0",x"E0",x"C0",x"00", -- 0x0510
		x"60",x"00",x"C0",x"00",x"F0",x"E0",x"70",x"E0", -- 0x0518
		x"00",x"00",x"C0",x"20",x"60",x"60",x"30",x"C0", -- 0x0520
		x"10",x"80",x"30",x"C0",x"60",x"60",x"C0",x"20", -- 0x0528
		x"00",x"00",x"00",x"E0",x"10",x"E0",x"F0",x"00", -- 0x0530
		x"F0",x"00",x"10",x"E0",x"00",x"E0",x"00",x"00", -- 0x0538
		x"00",x"00",x"80",x"20",x"C0",x"20",x"E0",x"20", -- 0x0540
		x"B0",x"20",x"90",x"A0",x"80",x"E0",x"80",x"60", -- 0x0548
		x"00",x"F0",x"10",x"00",x"00",x"C0",x"10",x"00", -- 0x0550
		x"90",x"F0",x"D0",x"00",x"B0",x"00",x"90",x"00", -- 0x0558
		x"10",x"10",x"00",x"B0",x"00",x"40",x"00",x"A0", -- 0x0560
		x"90",x"10",x"D0",x"10",x"B0",x"00",x"90",x"00", -- 0x0568
		x"00",x"30",x"00",x"40",x"30",x"80",x"00",x"40", -- 0x0570
		x"90",x"30",x"D0",x"00",x"B0",x"00",x"90",x"00", -- 0x0578
		x"00",x"F0",x"10",x"00",x"00",x"C0",x"10",x"00", -- 0x0580
		x"00",x"F0",x"30",x"00",x"C0",x"00",x"30",x"00", -- 0x0588
		x"20",x"10",x"10",x"30",x"00",x"C0",x"00",x"C0", -- 0x0590
		x"10",x"30",x"30",x"10",x"C0",x"00",x"30",x"00", -- 0x0598
		x"00",x"F0",x"10",x"00",x"00",x"C0",x"10",x"00", -- 0x05A0
		x"90",x"F0",x"60",x"00",x"60",x"00",x"90",x"00", -- 0x05A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40", -- 0x05B0
		x"00",x"30",x"00",x"30",x"00",x"00",x"00",x"00", -- 0x05B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05F8
		x"00",x"00",x"8F",x"0E",x"8F",x"0E",x"EF",x"CE", -- 0x0600
		x"23",x"46",x"23",x"0E",x"33",x"2E",x"11",x"CC", -- 0x0608
		x"00",x"00",x"11",x"FF",x"00",x"55",x"00",x"55", -- 0x0610
		x"0B",x"2A",x"0A",x"08",x"0A",x"08",x"04",x"00", -- 0x0618
		x"00",x"00",x"10",x"F0",x"1A",x"F0",x"0F",x"50", -- 0x0620
		x"08",x"50",x"06",x"70",x"09",x"20",x"06",x"00", -- 0x0628
		x"00",x"00",x"00",x"FF",x"01",x"55",x"0F",x"5D", -- 0x0630
		x"00",x"22",x"0B",x"08",x"0A",x"08",x"04",x"00", -- 0x0638
		x"00",x"00",x"09",x"F0",x"0C",x"58",x"0A",x"58", -- 0x0640
		x"09",x"20",x"07",x"00",x"08",x"08",x"07",x"00", -- 0x0648
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0650
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0658
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0660
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0668
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0670
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0678
		x"F8",x"F0",x"F8",x"F0",x"FF",x"F6",x"11",x"B2", -- 0x0680
		x"10",x"B2",x"F8",x"F0",x"F9",x"F9",x"EE",x"EE", -- 0x0688
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0690
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0698
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0700
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0708
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0710
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0718
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0720
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0728
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0730
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0738
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0740
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0748
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0750
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0760
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0768
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0770
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0798
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F8
		x"00",x"00",x"33",x"FF",x"33",x"FF",x"F3",x"FF", -- 0x0800
		x"F3",x"FF",x"F3",x"F0",x"F3",x"F0",x"F3",x"00", -- 0x0808
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0810
		x"FF",x"FF",x"F0",x"F3",x"F0",x"F3",x"00",x"F3", -- 0x0818
		x"F3",x"00",x"F3",x"00",x"F3",x"FF",x"F3",x"FF", -- 0x0820
		x"F3",x"FF",x"F3",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x0828
		x"00",x"F3",x"00",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x0830
		x"FF",x"FF",x"FF",x"FF",x"F0",x"C0",x"F0",x"C0", -- 0x0838
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0840
		x"00",x"00",x"00",x"00",x"00",x"00",x"33",x"FF", -- 0x0848
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0850
		x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF", -- 0x0858
		x"33",x"FF",x"F3",x"FF",x"F3",x"FF",x"F0",x"F0", -- 0x0860
		x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0868
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"C0", -- 0x0870
		x"F0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0878
		x"00",x"00",x"33",x"FF",x"33",x"FF",x"F3",x"FF", -- 0x0880
		x"F3",x"FF",x"F3",x"F0",x"F3",x"F0",x"F3",x"30", -- 0x0888
		x"00",x"00",x"CC",x"33",x"CC",x"33",x"CC",x"F3", -- 0x0890
		x"CC",x"F3",x"CC",x"F3",x"CC",x"F3",x"CC",x"F3", -- 0x0898
		x"F3",x"30",x"F3",x"30",x"F3",x"30",x"F3",x"30", -- 0x08A0
		x"F3",x"30",x"F3",x"30",x"C0",x"30",x"C0",x"30", -- 0x08A8
		x"CC",x"F3",x"CC",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x08B0
		x"FF",x"FF",x"FF",x"FF",x"F0",x"C0",x"F0",x"C0", -- 0x08B8
		x"00",x"00",x"33",x"00",x"33",x"00",x"F3",x"30", -- 0x08C0
		x"F3",x"30",x"F3",x"30",x"F3",x"30",x"F3",x"30", -- 0x08C8
		x"00",x"00",x"CC",x"33",x"CC",x"33",x"CC",x"F3", -- 0x08D0
		x"CC",x"F3",x"CC",x"F3",x"CC",x"F3",x"CC",x"F3", -- 0x08D8
		x"F3",x"30",x"F3",x"30",x"F3",x"FF",x"F3",x"FF", -- 0x08E0
		x"F3",x"FF",x"F3",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x08E8
		x"CC",x"F3",x"CC",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x08F0
		x"FF",x"FF",x"FF",x"FF",x"F0",x"C0",x"F0",x"C0", -- 0x08F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30", -- 0x0900
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x0908
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0910
		x"FF",x"FF",x"FC",x"C0",x"FC",x"C0",x"CC",x"00", -- 0x0918
		x"00",x"30",x"00",x"30",x"33",x"FF",x"33",x"FF", -- 0x0920
		x"F3",x"FF",x"F3",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x0928
		x"CC",x"00",x"CC",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x0930
		x"FF",x"FF",x"FF",x"FF",x"F0",x"C0",x"F0",x"C0", -- 0x0938
		x"00",x"00",x"33",x"00",x"33",x"00",x"F3",x"30", -- 0x0940
		x"F3",x"30",x"F3",x"30",x"F3",x"30",x"F3",x"30", -- 0x0948
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0950
		x"FF",x"FF",x"FC",x"F3",x"FC",x"F3",x"CC",x"F3", -- 0x0958
		x"F3",x"30",x"F3",x"30",x"F3",x"FF",x"F3",x"FF", -- 0x0960
		x"F3",x"FF",x"F3",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x0968
		x"CC",x"F3",x"CC",x"F3",x"CC",x"F3",x"CC",x"F3", -- 0x0970
		x"CC",x"F3",x"CC",x"F3",x"00",x"C0",x"00",x"C0", -- 0x0978
		x"00",x"00",x"33",x"FF",x"33",x"FF",x"F3",x"FF", -- 0x0980
		x"F3",x"FF",x"F3",x"F0",x"F3",x"F0",x"F3",x"30", -- 0x0988
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0990
		x"FF",x"FF",x"FC",x"F3",x"FC",x"F3",x"CC",x"F3", -- 0x0998
		x"F3",x"30",x"F3",x"30",x"F3",x"FF",x"F3",x"FF", -- 0x09A0
		x"F3",x"FF",x"F3",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x09A8
		x"CC",x"F3",x"CC",x"F3",x"CC",x"F3",x"CC",x"F3", -- 0x09B0
		x"CC",x"F3",x"CC",x"F3",x"00",x"C0",x"00",x"C0", -- 0x09B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09C8
		x"00",x"00",x"00",x"33",x"00",x"33",x"00",x"F3", -- 0x09D0
		x"00",x"F3",x"00",x"F3",x"00",x"F3",x"00",x"F3", -- 0x09D8
		x"00",x"00",x"00",x"00",x"33",x"FF",x"33",x"FF", -- 0x09E0
		x"F3",x"FF",x"F3",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x09E8
		x"00",x"F3",x"00",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x09F0
		x"FF",x"FF",x"FF",x"FF",x"F0",x"C0",x"F0",x"C0", -- 0x09F8
		x"00",x"00",x"33",x"FF",x"33",x"FF",x"F3",x"FF", -- 0x0A00
		x"F3",x"FF",x"F3",x"F0",x"F3",x"F0",x"F3",x"30", -- 0x0A08
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A10
		x"FF",x"FF",x"FC",x"F3",x"FC",x"F3",x"CC",x"F3", -- 0x0A18
		x"F3",x"30",x"F3",x"30",x"F3",x"FF",x"F3",x"FF", -- 0x0A20
		x"F3",x"FF",x"F3",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x0A28
		x"CC",x"F3",x"CC",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x0A30
		x"FF",x"FF",x"FF",x"FF",x"F0",x"C0",x"F0",x"C0", -- 0x0A38
		x"00",x"00",x"33",x"00",x"33",x"00",x"F3",x"30", -- 0x0A40
		x"F3",x"30",x"F3",x"30",x"F3",x"30",x"F3",x"30", -- 0x0A48
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A50
		x"FF",x"FF",x"FC",x"F3",x"FC",x"F3",x"CC",x"F3", -- 0x0A58
		x"F3",x"30",x"F3",x"30",x"F3",x"FF",x"F3",x"FF", -- 0x0A60
		x"F3",x"FF",x"F3",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x0A68
		x"CC",x"F3",x"CC",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x0A70
		x"FF",x"FF",x"FF",x"FF",x"F0",x"C0",x"F0",x"C0", -- 0x0A78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0AF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0B98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0ED0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0ED8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0F98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0FF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1000
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"08", -- 0x1008
		x"03",x"0F",x"03",x"0F",x"03",x"0F",x"03",x"0F", -- 0x1010
		x"03",x"0F",x"03",x"0F",x"03",x"1E",x"03",x"1E", -- 0x1018
		x"0F",x"00",x"0F",x"00",x"0F",x"00",x"0F",x"00", -- 0x1020
		x"0F",x"00",x"0F",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x1028
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1030
		x"00",x"00",x"00",x"00",x"87",x"0F",x"87",x"0F", -- 0x1038
		x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"07", -- 0x1040
		x"00",x"07",x"00",x"03",x"0F",x"0F",x"0F",x"0F", -- 0x1048
		x"03",x"0C",x"0F",x"0E",x"0F",x"0F",x"0F",x"0F", -- 0x1050
		x"0F",x"0F",x"0F",x"0F",x"0F",x"1E",x"0F",x"78", -- 0x1058
		x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00", -- 0x1060
		x"0C",x"00",x"48",x"00",x"E0",x"00",x"FC",x"00", -- 0x1068
		x"03",x"1E",x"03",x"1E",x"03",x"1E",x"03",x"1E", -- 0x1070
		x"03",x"1E",x"03",x"1E",x"03",x"1E",x"03",x"1E", -- 0x1078
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1080
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1088
		x"87",x"0F",x"87",x"0F",x"87",x"0F",x"87",x"0F", -- 0x1090
		x"87",x"0F",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x1098
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x10A0
		x"0F",x"0F",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x10A8
		x"1E",x"F3",x"78",x"F7",x"3C",x"FF",x"1E",x"FF", -- 0x10B0
		x"1E",x"F7",x"F0",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x10B8
		x"DC",x"80",x"CC",x"C0",x"CC",x"60",x"CC",x"20", -- 0x10C0
		x"CC",x"20",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x10C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10D0
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"FF",x"00", -- 0x10D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x10E8
		x"CC",x"20",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x10F0
		x"00",x"20",x"00",x"20",x"00",x"20",x"00",x"20", -- 0x10F8
		x"03",x"1E",x"03",x"1E",x"00",x"10",x"00",x"10", -- 0x1100
		x"00",x"10",x"00",x"10",x"00",x"10",x"00",x"10", -- 0x1108
		x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",x"00", -- 0x1110
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x1118
		x"F0",x"F0",x"F0",x"F0",x"80",x"00",x"80",x"00", -- 0x1120
		x"80",x"00",x"80",x"00",x"80",x"00",x"80",x"00", -- 0x1128
		x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00", -- 0x1130
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1138
		x"F0",x"E0",x"F0",x"E0",x"00",x"00",x"00",x"00", -- 0x1140
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1148
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1150
		x"00",x"00",x"00",x"00",x"03",x"0F",x"03",x"0F", -- 0x1158
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1160
		x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F", -- 0x1168
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1170
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01", -- 0x1178
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1180
		x"00",x"00",x"00",x"00",x"0F",x"00",x"0F",x"08", -- 0x1188
		x"03",x"0F",x"03",x"0F",x"03",x"0F",x"03",x"0F", -- 0x1190
		x"03",x"1E",x"03",x"1E",x"03",x"1E",x"03",x"1E", -- 0x1198
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x11A0
		x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x11A8
		x"00",x"03",x"00",x"07",x"00",x"0F",x"01",x"0F", -- 0x11B0
		x"F0",x"87",x"F0",x"87",x"33",x"87",x"33",x"87", -- 0x11B8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x11C0
		x"0F",x"78",x"0F",x"F3",x"1E",x"F7",x"3C",x"FF", -- 0x11C8
		x"0F",x"0C",x"0F",x"0E",x"0F",x"0F",x"0F",x"0F", -- 0x11D0
		x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00", -- 0x11E0
		x"80",x"00",x"C0",x"00",x"E8",x"00",x"FC",x"00", -- 0x11E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11F0
		x"FF",x"FF",x"FF",x"88",x"FF",x"88",x"FF",x"88", -- 0x11F8
		x"33",x"87",x"33",x"87",x"33",x"96",x"33",x"96", -- 0x1200
		x"33",x"96",x"33",x"96",x"33",x"96",x"33",x"96", -- 0x1208
		x"79",x"FF",x"F3",x"FF",x"F7",x"FF",x"FF",x"FF", -- 0x1210
		x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00", -- 0x1218
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1220
		x"FF",x"FF",x"77",x"FF",x"77",x"FF",x"77",x"FF", -- 0x1228
		x"DC",x"80",x"CC",x"C0",x"CC",x"60",x"CC",x"20", -- 0x1230
		x"CC",x"20",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x1238
		x"FF",x"88",x"FF",x"88",x"FF",x"88",x"FF",x"FF", -- 0x1240
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1248
		x"33",x"96",x"F0",x"96",x"F0",x"96",x"87",x"1E", -- 0x1250
		x"87",x"1E",x"87",x"1E",x"87",x"1E",x"87",x"1E", -- 0x1258
		x"FF",x"00",x"FF",x"00",x"FF",x"00",x"FF",x"FF", -- 0x1260
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1268
		x"77",x"FF",x"F0",x"F1",x"F7",x"FD",x"F7",x"FD", -- 0x1270
		x"F7",x"FD",x"F7",x"FD",x"F7",x"FD",x"F7",x"FD", -- 0x1278
		x"CC",x"20",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x1280
		x"CC",x"20",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x1288
		x"03",x"1E",x"03",x"1E",x"03",x"1E",x"03",x"1E", -- 0x1290
		x"01",x"1E",x"00",x"1E",x"00",x"16",x"00",x"12", -- 0x1298
		x"87",x"1E",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x12A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12A8
		x"F7",x"FD",x"F0",x"F1",x"FF",x"FF",x"FF",x"FF", -- 0x12B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"CC", -- 0x12B8
		x"CC",x"20",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x12C0
		x"88",x"20",x"00",x"20",x"00",x"20",x"00",x"20", -- 0x12C8
		x"00",x"10",x"00",x"10",x"00",x"00",x"00",x"00", -- 0x12D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12D8
		x"FF",x"FF",x"F7",x"FF",x"C0",x"00",x"60",x"00", -- 0x12E0
		x"30",x"00",x"10",x"80",x"00",x"F0",x"00",x"70", -- 0x12E8
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x12F0
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x12F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1300
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1308
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1310
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1318
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1320
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1328
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1330
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1338
		x"FF",x"88",x"FF",x"00",x"00",x"00",x"00",x"00", -- 0x1340
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x1348
		x"00",x"20",x"00",x"60",x"00",x"C0",x"10",x"80", -- 0x1350
		x"30",x"00",x"60",x"00",x"C0",x"00",x"80",x"00", -- 0x1358
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1360
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"01", -- 0x1368
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1370
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x1378
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1380
		x"00",x"00",x"0C",x"00",x"0E",x"00",x"0F",x"08", -- 0x1388
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"01", -- 0x1390
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"01", -- 0x1398
		x"0F",x"0F",x"0F",x"0F",x"1E",x"F0",x"1E",x"FF", -- 0x13A0
		x"1E",x"FF",x"1E",x"FF",x"1E",x"FF",x"1E",x"FF", -- 0x13A8
		x"0F",x"0E",x"0F",x"0F",x"F0",x"87",x"FF",x"E1", -- 0x13B0
		x"FF",x"F8",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x13B8
		x"00",x"00",x"00",x"00",x"0C",x"00",x"0E",x"00", -- 0x13C0
		x"87",x"00",x"C3",x"0C",x"F8",x"0F",x"FE",x"87", -- 0x13C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00", -- 0x13D8
		x"00",x"00",x"00",x"00",x"03",x"0F",x"03",x"0F", -- 0x13E0
		x"03",x"0F",x"03",x"0F",x"03",x"0F",x"03",x"0F", -- 0x13E8
		x"00",x"01",x"00",x"01",x"0F",x"01",x"0F",x"01", -- 0x13F0
		x"0F",x"01",x"0F",x"01",x"0F",x"01",x"0F",x"0F", -- 0x13F8
		x"1E",x"FF",x"1E",x"BB",x"1E",x"99",x"1E",x"88", -- 0x1400
		x"1E",x"88",x"1E",x"88",x"1E",x"88",x"1E",x"FF", -- 0x1408
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x1410
		x"33",x"FF",x"00",x"FF",x"60",x"77",x"F8",x"F7", -- 0x1418
		x"FF",x"E1",x"FF",x"FC",x"FF",x"FE",x"FF",x"FF", -- 0x1420
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1428
		x"0C",x"00",x"84",x"00",x"C0",x"00",x"F8",x"00", -- 0x1430
		x"DC",x"C0",x"CC",x"60",x"CC",x"20",x"CC",x"20", -- 0x1438
		x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x1440
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1448
		x"96",x"FF",x"96",x"FF",x"96",x"FF",x"96",x"FF", -- 0x1450
		x"96",x"FF",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1458
		x"FB",x"F1",x"FB",x"FC",x"FB",x"FE",x"FB",x"FF", -- 0x1460
		x"FB",x"FF",x"F8",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x1468
		x"FF",x"FF",x"FF",x"FF",x"F3",x"FF",x"F8",x"FF", -- 0x1470
		x"FE",x"F3",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x1478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1480
		x"FF",x"FF",x"FF",x"FF",x"FF",x"11",x"FF",x"11", -- 0x1488
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1490
		x"FF",x"FF",x"FF",x"FF",x"FF",x"88",x"FF",x"88", -- 0x1498
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14A0
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x14A8
		x"CC",x"20",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x14B0
		x"CC",x"20",x"CC",x"20",x"00",x"20",x"00",x"20", -- 0x14B8
		x"03",x"1E",x"03",x"1E",x"03",x"1E",x"00",x"10", -- 0x14C0
		x"00",x"10",x"00",x"10",x"00",x"10",x"00",x"10", -- 0x14C8
		x"FF",x"11",x"FF",x"11",x"FF",x"11",x"00",x"00", -- 0x14D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14D8
		x"FF",x"88",x"FF",x"88",x"FF",x"88",x"F0",x"00", -- 0x14E0
		x"90",x"00",x"90",x"00",x"90",x"00",x"90",x"00", -- 0x14E8
		x"00",x"00",x"00",x"00",x"70",x"F0",x"70",x"F0", -- 0x14F0
		x"40",x"00",x"40",x"00",x"40",x"00",x"40",x"00", -- 0x14F8
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x1500
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1508
		x"00",x"20",x"00",x"20",x"F0",x"E0",x"F0",x"E0", -- 0x1510
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1518
		x"00",x"10",x"00",x"10",x"00",x"00",x"00",x"00", -- 0x1520
		x"00",x"00",x"03",x"0F",x"03",x"0F",x"03",x"0F", -- 0x1528
		x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00", -- 0x1530
		x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x1538
		x"90",x"F0",x"90",x"F0",x"00",x"00",x"00",x"00", -- 0x1540
		x"00",x"00",x"0F",x"00",x"0F",x"00",x"0F",x"08", -- 0x1548
		x"C0",x"00",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x1550
		x"00",x"00",x"00",x"0F",x"00",x"0F",x"00",x"0F", -- 0x1558
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1560
		x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x1568
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1570
		x"00",x"00",x"0C",x"00",x"0C",x"00",x"0C",x"00", -- 0x1578
		x"03",x"0F",x"03",x"0F",x"03",x"0F",x"03",x"1E", -- 0x1580
		x"03",x"1E",x"03",x"1E",x"03",x"1E",x"03",x"1E", -- 0x1588
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0", -- 0x1590
		x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1598
		x"0F",x"08",x"0F",x"08",x"0F",x"0C",x"F0",x"F0", -- 0x15A0
		x"F0",x"F0",x"FF",x"FE",x"FF",x"EE",x"FF",x"EE", -- 0x15A8
		x"00",x"0F",x"00",x"0F",x"00",x"0F",x"00",x"0F", -- 0x15B0
		x"00",x"0F",x"80",x"0F",x"80",x"0F",x"C0",x"0F", -- 0x15B8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0", -- 0x15C0
		x"F0",x"F0",x"F7",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x15C8
		x"0C",x"00",x"0C",x"00",x"0C",x"00",x"F0",x"E0", -- 0x15D0
		x"F0",x"E0",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x15D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"99", -- 0x15E0
		x"FF",x"99",x"FF",x"88",x"FF",x"88",x"FF",x"88", -- 0x15E8
		x"40",x"0F",x"40",x"0F",x"E8",x"0F",x"A8",x"00", -- 0x15F0
		x"B8",x"00",x"DC",x"00",x"DC",x"00",x"FE",x"80", -- 0x15F8
		x"F7",x"FF",x"F7",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x1600
		x"F7",x"FF",x"F7",x"FF",x"F7",x"FF",x"F0",x"F3", -- 0x1608
		x"FF",x"88",x"FF",x"88",x"FF",x"88",x"FF",x"FF", -- 0x1610
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1618
		x"F0",x"FF",x"96",x"F7",x"83",x"F7",x"83",x"F3", -- 0x1620
		x"81",x"7B",x"81",x"79",x"81",x"3D",x"80",x"3C", -- 0x1628
		x"EE",x"80",x"EE",x"C0",x"FF",x"40",x"FF",x"CB", -- 0x1630
		x"FF",x"E9",x"FF",x"ED",x"FF",x"FC",x"FF",x"FE", -- 0x1638
		x"F0",x"F3",x"0F",x"7B",x"0F",x"7B",x"0F",x"7B", -- 0x1640
		x"0F",x"7B",x"0F",x"7B",x"0F",x"7B",x"0F",x"7B", -- 0x1648
		x"80",x"1E",x"F0",x"96",x"88",x"96",x"88",x"83", -- 0x1650
		x"88",x"83",x"88",x"83",x"88",x"81",x"88",x"81", -- 0x1658
		x"FF",x"FE",x"FF",x"FE",x"F7",x"FF",x"F7",x"FF", -- 0x1660
		x"F3",x"FF",x"7B",x"FF",x"79",x"FF",x"79",x"FF", -- 0x1668
		x"0F",x"7B",x"F0",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x1670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"CC", -- 0x1678
		x"CC",x"20",x"CC",x"20",x"CC",x"20",x"CC",x"20", -- 0x1680
		x"88",x"20",x"00",x"20",x"00",x"20",x"00",x"20", -- 0x1688
		x"03",x"1E",x"03",x"1E",x"00",x"10",x"00",x"10", -- 0x1690
		x"00",x"10",x"00",x"10",x"00",x"10",x"00",x"10", -- 0x1698
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x16A0
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x16A8
		x"88",x"80",x"88",x"80",x"00",x"80",x"00",x"80", -- 0x16B0
		x"00",x"80",x"00",x"80",x"F0",x"80",x"F0",x"80", -- 0x16B8
		x"3D",x"FF",x"30",x"00",x"10",x"00",x"10",x"80", -- 0x16C0
		x"00",x"80",x"00",x"C0",x"00",x"70",x"00",x"30", -- 0x16C8
		x"FF",x"88",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D0
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x16D8
		x"00",x"20",x"00",x"60",x"00",x"C0",x"10",x"80", -- 0x16E0
		x"30",x"00",x"60",x"00",x"C0",x"00",x"80",x"00", -- 0x16E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1700
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1708
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1710
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1718
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1720
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1728
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1730
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1738
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1740
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1748
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1750
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1760
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1768
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1770
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1778
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1798
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1800
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1808
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1810
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1818
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1820
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1828
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1830
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1838
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1840
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1848
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1850
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1858
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1860
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1868
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1870
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1878
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1880
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1888
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1890
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1898
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1900
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1908
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1910
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1918
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1920
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1928
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1930
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1938
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1940
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1948
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1950
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1958
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1960
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1968
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1970
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1978
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1980
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1988
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1990
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1998
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
		x"00",x"00",x"03",x"08",x"04",x"04",x"09",x"02", -- 0x1F90
		x"0A",x"0A",x"0A",x"0A",x"04",x"04",x"03",x"08", -- 0x1F98
		x"00",x"00",x"07",x"0C",x"0F",x"0E",x"08",x"02", -- 0x1FA0
		x"08",x"02",x"08",x"06",x"0C",x"04",x"04",x"00", -- 0x1FA8
		x"00",x"00",x"0F",x"08",x"0F",x"0C",x"02",x"06", -- 0x1FB0
		x"02",x"02",x"02",x"06",x"0F",x"0C",x"0F",x"08", -- 0x1FB8
		x"00",x"00",x"0F",x"0E",x"0F",x"0E",x"01",x"02", -- 0x1FC0
		x"01",x"02",x"01",x"02",x"01",x"0E",x"00",x"0C", -- 0x1FC8
		x"00",x"00",x"07",x"0C",x"0F",x"0E",x"08",x"02", -- 0x1FD0
		x"08",x"02",x"08",x"06",x"0C",x"04",x"04",x"00", -- 0x1FD8
		x"00",x"00",x"07",x"0C",x"0F",x"0E",x"08",x"02", -- 0x1FE0
		x"08",x"02",x"08",x"02",x"0F",x"0E",x"07",x"0C", -- 0x1FE8
		x"00",x"00",x"0F",x"0E",x"0F",x"0E",x"00",x"0C", -- 0x1FF0
		x"01",x"08",x"00",x"0C",x"0F",x"0E",x"0F",x"0E"  -- 0x1FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
