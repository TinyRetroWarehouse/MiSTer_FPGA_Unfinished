-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_M5 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_M5 is


	type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"84",x"B0",x"84",x"31",x"85",x"76",x"85",x"D3", -- 0x0000
		x"85",x"30",x"86",x"91",x"86",x"1E",x"28",x"00", -- 0x0008
		x"02",x"05",x"29",x"00",x"02",x"05",x"2A",x"00", -- 0x0010
		x"02",x"05",x"2B",x"00",x"02",x"05",x"2C",x"00", -- 0x0018
		x"02",x"05",x"2D",x"00",x"02",x"05",x"2E",x"00", -- 0x0020
		x"02",x"05",x"2F",x"00",x"02",x"0A",x"48",x"00", -- 0x0028
		x"02",x"01",x"49",x"00",x"02",x"02",x"49",x"00", -- 0x0030
		x"01",x"01",x"49",x"00",x"02",x"03",x"49",x"00", -- 0x0038
		x"01",x"01",x"49",x"FF",x"01",x"02",x"49",x"00", -- 0x0040
		x"01",x"02",x"49",x"FF",x"01",x"01",x"4A",x"FF", -- 0x0048
		x"01",x"01",x"4A",x"FF",x"00",x"01",x"4A",x"FF", -- 0x0050
		x"01",x"04",x"4A",x"FF",x"00",x"01",x"4A",x"FF", -- 0x0058
		x"FF",x"01",x"4B",x"FF",x"00",x"03",x"4B",x"FF", -- 0x0060
		x"FF",x"02",x"4B",x"00",x"FF",x"01",x"4B",x"FF", -- 0x0068
		x"FF",x"02",x"4C",x"00",x"FF",x"01",x"4C",x"00", -- 0x0070
		x"FE",x"02",x"4C",x"00",x"FF",x"13",x"1C",x"00", -- 0x0078
		x"FE",x"05",x"1D",x"00",x"FE",x"05",x"1E",x"00", -- 0x0080
		x"FE",x"05",x"1F",x"00",x"FE",x"05",x"18",x"00", -- 0x0088
		x"FE",x"05",x"19",x"00",x"FE",x"05",x"1A",x"00", -- 0x0090
		x"FE",x"05",x"1B",x"00",x"FE",x"04",x"1C",x"00", -- 0x0098
		x"FE",x"01",x"4C",x"00",x"FE",x"02",x"4C",x"00", -- 0x00A0
		x"FF",x"01",x"4C",x"00",x"FE",x"03",x"4C",x"00", -- 0x00A8
		x"FF",x"01",x"4C",x"FF",x"FF",x"02",x"4C",x"00", -- 0x00B0
		x"FF",x"02",x"4C",x"FF",x"FF",x"01",x"4B",x"FF", -- 0x00B8
		x"FF",x"01",x"4B",x"FF",x"00",x"01",x"4B",x"FF", -- 0x00C0
		x"FF",x"04",x"4B",x"FF",x"00",x"01",x"4B",x"FF", -- 0x00C8
		x"FF",x"01",x"4A",x"FF",x"00",x"03",x"4A",x"FF", -- 0x00D0
		x"01",x"02",x"4A",x"00",x"01",x"01",x"4A",x"FF", -- 0x00D8
		x"01",x"02",x"49",x"00",x"01",x"01",x"49",x"00", -- 0x00E0
		x"02",x"02",x"49",x"00",x"01",x"17",x"28",x"00", -- 0x00E8
		x"02",x"05",x"29",x"00",x"02",x"05",x"2A",x"00", -- 0x00F0
		x"02",x"05",x"2B",x"00",x"02",x"05",x"2C",x"00", -- 0x00F8
		x"02",x"05",x"2D",x"00",x"02",x"05",x"2E",x"00", -- 0x0100
		x"02",x"05",x"2F",x"00",x"02",x"63",x"28",x"00", -- 0x0108
		x"02",x"00",x"18",x"0C",x"00",x"02",x"01",x"0B", -- 0x0110
		x"FF",x"03",x"01",x"0B",x"00",x"02",x"03",x"0B", -- 0x0118
		x"FF",x"03",x"02",x"0B",x"FF",x"02",x"01",x"0A", -- 0x0120
		x"FE",x"02",x"01",x"0A",x"FF",x"02",x"03",x"0A", -- 0x0128
		x"FE",x"02",x"01",x"09",x"FD",x"01",x"02",x"09", -- 0x0130
		x"FE",x"01",x"01",x"09",x"FD",x"01",x"01",x"09", -- 0x0138
		x"FE",x"01",x"04",x"08",x"FE",x"00",x"01",x"07", -- 0x0140
		x"FE",x"FF",x"01",x"07",x"FD",x"FF",x"02",x"07", -- 0x0148
		x"FE",x"FF",x"01",x"07",x"FD",x"FF",x"03",x"06", -- 0x0150
		x"FE",x"FE",x"01",x"06",x"FF",x"FE",x"01",x"06", -- 0x0158
		x"FE",x"FE",x"02",x"05",x"FF",x"FE",x"03",x"05", -- 0x0160
		x"FF",x"FD",x"01",x"05",x"00",x"FE",x"01",x"05", -- 0x0168
		x"FF",x"FD",x"08",x"04",x"00",x"FE",x"01",x"03", -- 0x0170
		x"01",x"FD",x"01",x"03",x"00",x"FE",x"03",x"03", -- 0x0178
		x"01",x"FD",x"02",x"03",x"01",x"FE",x"01",x"02", -- 0x0180
		x"02",x"FE",x"01",x"02",x"01",x"FE",x"03",x"02", -- 0x0188
		x"02",x"FE",x"01",x"01",x"03",x"FF",x"02",x"01", -- 0x0190
		x"02",x"FF",x"01",x"01",x"03",x"FF",x"01",x"01", -- 0x0198
		x"02",x"FF",x"04",x"00",x"02",x"00",x"01",x"0F", -- 0x01A0
		x"02",x"01",x"01",x"0F",x"03",x"01",x"02",x"0F", -- 0x01A8
		x"02",x"01",x"01",x"0F",x"03",x"01",x"03",x"0E", -- 0x01B0
		x"02",x"02",x"01",x"0E",x"01",x"02",x"01",x"0E", -- 0x01B8
		x"02",x"02",x"02",x"0D",x"01",x"02",x"03",x"0D", -- 0x01C0
		x"01",x"03",x"01",x"0D",x"00",x"02",x"01",x"0D", -- 0x01C8
		x"01",x"03",x"04",x"0C",x"00",x"02",x"3C",x"0C", -- 0x01D0
		x"00",x"02",x"01",x"0B",x"FF",x"03",x"01",x"0B", -- 0x01D8
		x"00",x"02",x"03",x"0B",x"FF",x"03",x"02",x"0B", -- 0x01E0
		x"FF",x"02",x"01",x"0A",x"FE",x"02",x"01",x"0A", -- 0x01E8
		x"FF",x"02",x"03",x"0A",x"FE",x"02",x"01",x"09", -- 0x01F0
		x"FD",x"01",x"02",x"09",x"FE",x"01",x"01",x"09", -- 0x01F8
		x"FD",x"01",x"01",x"09",x"FE",x"01",x"04",x"08", -- 0x0200
		x"FE",x"00",x"01",x"07",x"FE",x"FF",x"01",x"07", -- 0x0208
		x"FD",x"FF",x"02",x"07",x"FE",x"FF",x"01",x"07", -- 0x0210
		x"FD",x"FF",x"03",x"06",x"FE",x"FE",x"01",x"06", -- 0x0218
		x"FF",x"FE",x"01",x"06",x"FE",x"FE",x"02",x"05", -- 0x0220
		x"FF",x"FE",x"03",x"05",x"FF",x"FD",x"01",x"05", -- 0x0228
		x"00",x"FE",x"01",x"05",x"FF",x"FD",x"08",x"04", -- 0x0230
		x"00",x"FE",x"01",x"03",x"01",x"FD",x"01",x"03", -- 0x0238
		x"00",x"FE",x"03",x"03",x"01",x"FD",x"02",x"03", -- 0x0240
		x"01",x"FE",x"01",x"02",x"02",x"FE",x"01",x"02", -- 0x0248
		x"01",x"FE",x"03",x"02",x"02",x"FE",x"01",x"01", -- 0x0250
		x"03",x"FF",x"02",x"01",x"02",x"FF",x"01",x"01", -- 0x0258
		x"03",x"FF",x"01",x"01",x"02",x"FF",x"04",x"00", -- 0x0260
		x"02",x"00",x"01",x"0F",x"02",x"01",x"01",x"0F", -- 0x0268
		x"03",x"01",x"02",x"0F",x"02",x"01",x"01",x"0F", -- 0x0270
		x"03",x"01",x"03",x"0E",x"02",x"02",x"01",x"0E", -- 0x0278
		x"01",x"02",x"01",x"0E",x"02",x"02",x"02",x"0D", -- 0x0280
		x"01",x"02",x"03",x"0D",x"01",x"03",x"01",x"0D", -- 0x0288
		x"00",x"02",x"01",x"0D",x"01",x"03",x"04",x"0C", -- 0x0290
		x"00",x"02",x"63",x"0C",x"00",x"02",x"00",x"37", -- 0x0298
		x"48",x"00",x"02",x"06",x"49",x"00",x"02",x"04", -- 0x02A0
		x"4A",x"00",x"02",x"04",x"4A",x"00",x"01",x"05", -- 0x02A8
		x"4A",x"00",x"00",x"04",x"4A",x"00",x"FF",x"04", -- 0x02B0
		x"4A",x"00",x"FE",x"06",x"4B",x"00",x"FE",x"19", -- 0x02B8
		x"4C",x"00",x"FE",x"06",x"4D",x"00",x"FE",x"04", -- 0x02C0
		x"4E",x"00",x"FE",x"04",x"4E",x"00",x"FF",x"04", -- 0x02C8
		x"4E",x"00",x"00",x"04",x"4E",x"00",x"01",x"04", -- 0x02D0
		x"4E",x"00",x"02",x"06",x"4F",x"00",x"02",x"63", -- 0x02D8
		x"48",x"00",x"02",x"00",x"28",x"48",x"00",x"02", -- 0x02E0
		x"02",x"49",x"00",x"01",x"02",x"49",x"00",x"00", -- 0x02E8
		x"02",x"4A",x"00",x"00",x"02",x"4A",x"00",x"FF", -- 0x02F0
		x"02",x"4A",x"00",x"FE",x"04",x"4B",x"00",x"FE", -- 0x02F8
		x"1E",x"4C",x"00",x"FE",x"04",x"4D",x"00",x"FE", -- 0x0300
		x"02",x"4E",x"00",x"FE",x"02",x"4E",x"00",x"FF", -- 0x0308
		x"02",x"4E",x"00",x"00",x"02",x"4F",x"00",x"00", -- 0x0310
		x"02",x"4F",x"00",x"01",x"06",x"4F",x"00",x"02", -- 0x0318
		x"63",x"48",x"00",x"02",x"00",x"22",x"0C",x"00", -- 0x0320
		x"02",x"01",x"0D",x"01",x"03",x"02",x"0D",x"00", -- 0x0328
		x"02",x"04",x"0D",x"01",x"03",x"04",x"0E",x"02", -- 0x0330
		x"02",x"04",x"0F",x"02",x"01",x"01",x"0F",x"03", -- 0x0338
		x"01",x"02",x"00",x"02",x"00",x"01",x"01",x"03", -- 0x0340
		x"FF",x"03",x"01",x"02",x"FE",x"02",x"02",x"01", -- 0x0348
		x"FE",x"04",x"02",x"01",x"FD",x"02",x"03",x"00", -- 0x0350
		x"FE",x"01",x"03",x"01",x"FD",x"05",x"04",x"00", -- 0x0358
		x"FE",x"01",x"05",x"FF",x"FE",x"02",x"05",x"00", -- 0x0360
		x"FE",x"03",x"05",x"FF",x"FE",x"01",x"06",x"FF", -- 0x0368
		x"FD",x"04",x"06",x"FE",x"FE",x"03",x"07",x"FE", -- 0x0370
		x"FF",x"02",x"07",x"FD",x"FF",x"01",x"07",x"FE", -- 0x0378
		x"FF",x"04",x"08",x"FE",x"00",x"04",x"09",x"FE", -- 0x0380
		x"01",x"06",x"0A",x"FE",x"02",x"03",x"0B",x"FF", -- 0x0388
		x"02",x"01",x"0B",x"FE",x"02",x"03",x"0B",x"FF", -- 0x0390
		x"02",x"03",x"0B",x"FF",x"03",x"01",x"0B",x"00", -- 0x0398
		x"02",x"02",x"0B",x"FF",x"03",x"04",x"0C",x"00", -- 0x03A0
		x"02",x"00",x"22",x"0C",x"00",x"02",x"01",x"0B", -- 0x03A8
		x"FF",x"03",x"02",x"0B",x"00",x"02",x"04",x"0B", -- 0x03B0
		x"FF",x"03",x"04",x"0A",x"FE",x"02",x"04",x"09", -- 0x03B8
		x"FE",x"01",x"01",x"09",x"FD",x"01",x"02",x"08", -- 0x03C0
		x"FE",x"00",x"01",x"07",x"FD",x"FF",x"03",x"07", -- 0x03C8
		x"FE",x"FE",x"02",x"06",x"FF",x"FE",x"04",x"06", -- 0x03D0
		x"FF",x"FD",x"02",x"05",x"00",x"FE",x"01",x"05", -- 0x03D8
		x"FF",x"FD",x"05",x"04",x"00",x"FE",x"01",x"03", -- 0x03E0
		x"01",x"FE",x"02",x"03",x"00",x"FE",x"03",x"03", -- 0x03E8
		x"01",x"FE",x"01",x"02",x"01",x"FD",x"04",x"02", -- 0x03F0
		x"02",x"FE",x"03",x"01",x"02",x"FF",x"02",x"01", -- 0x03F8
		x"03",x"FF",x"01",x"01",x"02",x"FF",x"04",x"00", -- 0x0400
		x"02",x"00",x"04",x"0F",x"02",x"01",x"06",x"0E", -- 0x0408
		x"02",x"02",x"03",x"0D",x"01",x"02",x"01",x"0D", -- 0x0410
		x"02",x"02",x"03",x"0D",x"01",x"02",x"03",x"0D", -- 0x0418
		x"01",x"03",x"01",x"0D",x"00",x"02",x"02",x"0D", -- 0x0420
		x"01",x"03",x"04",x"0C",x"00",x"02",x"00",x"22", -- 0x0428
		x"0C",x"00",x"02",x"01",x"0D",x"01",x"03",x"02", -- 0x0430
		x"0D",x"00",x"02",x"04",x"0D",x"01",x"03",x"04", -- 0x0438
		x"0E",x"02",x"02",x"04",x"0F",x"02",x"01",x"01", -- 0x0440
		x"0F",x"03",x"01",x"02",x"00",x"02",x"00",x"01", -- 0x0448
		x"01",x"03",x"FF",x"03",x"01",x"02",x"FE",x"02", -- 0x0450
		x"02",x"01",x"FE",x"04",x"02",x"01",x"FD",x"02", -- 0x0458
		x"03",x"00",x"FE",x"01",x"03",x"01",x"FD",x"05", -- 0x0460
		x"04",x"00",x"FE",x"01",x"05",x"FF",x"FE",x"02", -- 0x0468
		x"05",x"00",x"FE",x"03",x"05",x"FF",x"FE",x"01", -- 0x0470
		x"06",x"FF",x"FD",x"04",x"06",x"FE",x"FE",x"03", -- 0x0478
		x"07",x"FE",x"FF",x"02",x"07",x"FD",x"FF",x"01", -- 0x0480
		x"07",x"FE",x"FF",x"06",x"08",x"FE",x"00",x"01", -- 0x0488
		x"09",x"FF",x"01",x"04",x"09",x"FE",x"01",x"05", -- 0x0490
		x"0A",x"FE",x"02",x"03",x"0A",x"FF",x"02",x"06", -- 0x0498
		x"0B",x"FF",x"03",x"01",x"0B",x"00",x"02",x"01", -- 0x04A0
		x"0B",x"FF",x"03",x"06",x"0C",x"00",x"02",x"00", -- 0x04A8
		x"22",x"0C",x"00",x"02",x"01",x"0B",x"FF",x"03", -- 0x04B0
		x"02",x"0B",x"00",x"02",x"04",x"0B",x"FF",x"03", -- 0x04B8
		x"04",x"0A",x"FE",x"02",x"04",x"09",x"FE",x"01", -- 0x04C0
		x"01",x"09",x"FD",x"01",x"02",x"08",x"FE",x"00", -- 0x04C8
		x"01",x"07",x"FD",x"FF",x"03",x"07",x"FE",x"FE", -- 0x04D0
		x"02",x"06",x"FF",x"FE",x"04",x"06",x"FF",x"FD", -- 0x04D8
		x"02",x"05",x"00",x"FE",x"01",x"05",x"FF",x"FD", -- 0x04E0
		x"05",x"04",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x04E8
		x"02",x"03",x"00",x"FE",x"03",x"03",x"01",x"FE", -- 0x04F0
		x"01",x"02",x"01",x"FD",x"04",x"02",x"02",x"FE", -- 0x04F8
		x"03",x"01",x"02",x"FF",x"02",x"01",x"03",x"FF", -- 0x0500
		x"01",x"01",x"02",x"FF",x"06",x"00",x"02",x"00", -- 0x0508
		x"01",x"0F",x"01",x"01",x"04",x"0F",x"02",x"01", -- 0x0510
		x"05",x"0E",x"02",x"02",x"03",x"0E",x"01",x"02", -- 0x0518
		x"06",x"0D",x"01",x"03",x"01",x"0D",x"00",x"02", -- 0x0520
		x"01",x"0D",x"01",x"03",x"06",x"0C",x"00",x"02", -- 0x0528
		x"00",x"2C",x"40",x"FE",x"00",x"03",x"41",x"FE", -- 0x0530
		x"00",x"02",x"41",x"FF",x"00",x"02",x"41",x"00", -- 0x0538
		x"00",x"02",x"42",x"00",x"00",x"02",x"42",x"01", -- 0x0540
		x"00",x"03",x"42",x"02",x"00",x"03",x"43",x"02", -- 0x0548
		x"00",x"1C",x"44",x"02",x"00",x"03",x"45",x"03", -- 0x0550
		x"00",x"03",x"46",x"03",x"00",x"01",x"46",x"01", -- 0x0558
		x"00",x"02",x"46",x"00",x"00",x"02",x"47",x"00", -- 0x0560
		x"00",x"01",x"47",x"FF",x"00",x"03",x"47",x"FE", -- 0x0568
		x"00",x"63",x"40",x"FE",x"00",x"00",x"35",x"08", -- 0x0570
		x"FE",x"00",x"02",x"09",x"FE",x"01",x"03",x"0A", -- 0x0578
		x"FE",x"02",x"04",x"0B",x"FF",x"02",x"0C",x"0C", -- 0x0580
		x"00",x"02",x"02",x"0D",x"01",x"03",x"05",x"0E", -- 0x0588
		x"02",x"02",x"04",x"0F",x"03",x"01",x"0F",x"00", -- 0x0590
		x"02",x"00",x"02",x"01",x"03",x"FF",x"01",x"01", -- 0x0598
		x"02",x"FF",x"02",x"02",x"02",x"FE",x"04",x"03", -- 0x05A0
		x"01",x"FD",x"07",x"04",x"00",x"FE",x"04",x"05", -- 0x05A8
		x"FF",x"FE",x"02",x"06",x"FE",x"FE",x"03",x"07", -- 0x05B0
		x"FE",x"FF",x"08",x"08",x"FE",x"00",x"01",x"09", -- 0x05B8
		x"FD",x"01",x"04",x"09",x"FE",x"02",x"04",x"0A", -- 0x05C0
		x"FF",x"02",x"03",x"0B",x"FF",x"03",x"01",x"0C", -- 0x05C8
		x"00",x"02",x"00",x"35",x"08",x"FE",x"00",x"02", -- 0x05D0
		x"07",x"FE",x"FF",x"03",x"06",x"FE",x"FE",x"04", -- 0x05D8
		x"05",x"FF",x"FE",x"0C",x"04",x"00",x"FE",x"02", -- 0x05E0
		x"03",x"01",x"FD",x"05",x"02",x"02",x"FE",x"04", -- 0x05E8
		x"01",x"03",x"FF",x"0F",x"00",x"02",x"00",x"02", -- 0x05F0
		x"0F",x"03",x"01",x"01",x"0F",x"02",x"01",x"02", -- 0x05F8
		x"0E",x"02",x"02",x"04",x"0D",x"01",x"03",x"07", -- 0x0600
		x"0C",x"00",x"02",x"04",x"0B",x"FF",x"02",x"02", -- 0x0608
		x"0A",x"FE",x"02",x"03",x"09",x"FE",x"01",x"08", -- 0x0610
		x"08",x"FE",x"00",x"01",x"07",x"FD",x"FF",x"04", -- 0x0618
		x"07",x"FE",x"FE",x"04",x"06",x"FF",x"FE",x"03", -- 0x0620
		x"05",x"FF",x"FD",x"01",x"04",x"00",x"FE",x"00", -- 0x0628
		x"2C",x"08",x"FE",x"00",x"02",x"09",x"FD",x"01", -- 0x0630
		x"03",x"0A",x"FE",x"02",x"04",x"0B",x"FF",x"03", -- 0x0638
		x"0D",x"0C",x"00",x"02",x"04",x"0D",x"01",x"03", -- 0x0640
		x"05",x"0E",x"02",x"01",x"01",x"0F",x"03",x"01", -- 0x0648
		x"0D",x"00",x"02",x"00",x"02",x"01",x"02",x"FF", -- 0x0650
		x"03",x"02",x"02",x"FE",x"03",x"03",x"01",x"FD", -- 0x0658
		x"06",x"04",x"00",x"FE",x"03",x"05",x"FF",x"FD", -- 0x0660
		x"01",x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FE", -- 0x0668
		x"02",x"06",x"FE",x"FE",x"02",x"07",x"FE",x"FF", -- 0x0670
		x"04",x"08",x"FE",x"00",x"04",x"09",x"FE",x"01", -- 0x0678
		x"02",x"0A",x"FE",x"02",x"04",x"0B",x"FF",x"02", -- 0x0680
		x"02",x"0B",x"FF",x"03",x"01",x"0C",x"00",x"02", -- 0x0688
		x"00",x"2C",x"08",x"FE",x"00",x"02",x"07",x"FD", -- 0x0690
		x"FF",x"03",x"06",x"FE",x"FE",x"04",x"05",x"FF", -- 0x0698
		x"FD",x"0D",x"04",x"00",x"FE",x"04",x"03",x"01", -- 0x06A0
		x"FD",x"05",x"02",x"02",x"FF",x"01",x"01",x"03", -- 0x06A8
		x"FF",x"0D",x"00",x"02",x"00",x"02",x"0F",x"02", -- 0x06B0
		x"01",x"03",x"0E",x"02",x"02",x"03",x"0D",x"01", -- 0x06B8
		x"03",x"06",x"0C",x"00",x"02",x"03",x"0B",x"FF", -- 0x06C0
		x"03",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x06C8
		x"02",x"02",x"0A",x"FE",x"02",x"02",x"09",x"FE", -- 0x06D0
		x"01",x"04",x"08",x"FE",x"00",x"04",x"07",x"FE", -- 0x06D8
		x"FF",x"02",x"06",x"FE",x"FE",x"04",x"05",x"FF", -- 0x06E0
		x"FE",x"02",x"05",x"FF",x"FD",x"01",x"04",x"00", -- 0x06E8
		x"FE",x"00",x"FC",x"86",x"FC",x"86",x"10",x"87", -- 0x06F0
		x"24",x"87",x"38",x"87",x"00",x"00",x"00",x"04", -- 0x06F8
		x"00",x"00",x"10",x"04",x"00",x"00",x"20",x"04", -- 0x0700
		x"00",x"00",x"30",x"04",x"00",x"00",x"40",x"04", -- 0x0708
		x"00",x"00",x"00",x"04",x"10",x"00",x"10",x"04", -- 0x0710
		x"20",x"00",x"20",x"04",x"30",x"00",x"30",x"04", -- 0x0718
		x"40",x"00",x"40",x"04",x"00",x"00",x"00",x"04", -- 0x0720
		x"08",x"00",x"10",x"04",x"F8",x"00",x"10",x"04", -- 0x0728
		x"10",x"00",x"20",x"04",x"F0",x"00",x"20",x"04", -- 0x0730
		x"00",x"00",x"00",x"14",x"00",x"08",x"10",x"14", -- 0x0738
		x"00",x"F8",x"10",x"14",x"00",x"10",x"20",x"14", -- 0x0740
		x"00",x"F0",x"20",x"14",x"01",x"0E",x"01",x"0C", -- 0x0748
		x"01",x"0A",x"00",x"01",x"0A",x"01",x"09",x"01", -- 0x0750
		x"08",x"01",x"06",x"01",x"04",x"01",x"03",x"01", -- 0x0758
		x"02",x"01",x"01",x"01",x"00",x"00",x"04",x"00", -- 0x0760
		x"60",x"03",x"00",x"80",x"04",x"00",x"60",x"04", -- 0x0768
		x"08",x"40",x"04",x"08",x"20",x"02",x"08",x"00", -- 0x0770
		x"02",x"09",x"00",x"04",x"09",x"21",x"04",x"0A", -- 0x0778
		x"41",x"04",x"0A",x"61",x"FF",x"0B",x"81",x"03", -- 0x0780
		x"D8",x"05",x"D9",x"05",x"DA",x"05",x"DB",x"05", -- 0x0788
		x"DC",x"05",x"D9",x"05",x"DA",x"05",x"DB",x"05", -- 0x0790
		x"DC",x"05",x"DD",x"00",x"BA",x"87",x"BE",x"87", -- 0x0798
		x"C6",x"87",x"CE",x"87",x"D6",x"87",x"DE",x"87", -- 0x07A0
		x"BE",x"87",x"C2",x"87",x"C6",x"87",x"CA",x"87", -- 0x07A8
		x"CE",x"87",x"D2",x"87",x"D6",x"87",x"DA",x"87", -- 0x07B0
		x"DE",x"87",x"E2",x"87",x"1B",x"88",x"54",x"88", -- 0x07B8
		x"99",x"88",x"DE",x"88",x"53",x"89",x"C8",x"89", -- 0x07C0
		x"31",x"8A",x"9A",x"8A",x"07",x"8B",x"74",x"8B", -- 0x07C8
		x"E1",x"8B",x"4E",x"8C",x"C7",x"8C",x"40",x"8D", -- 0x07D0
		x"B1",x"8D",x"22",x"8E",x"A3",x"8E",x"24",x"8F", -- 0x07D8
		x"01",x"90",x"05",x"00",x"02",x"00",x"01",x"00", -- 0x07E0
		x"02",x"FF",x"01",x"01",x"02",x"00",x"05",x"01", -- 0x07E8
		x"02",x"FF",x"01",x"01",x"02",x"FE",x"01",x"02", -- 0x07F0
		x"02",x"FF",x"01",x"02",x"02",x"FE",x"01",x"02", -- 0x07F8
		x"01",x"FE",x"01",x"02",x"02",x"FE",x"01",x"02", -- 0x0800
		x"01",x"FE",x"05",x"03",x"01",x"FE",x"01",x"03", -- 0x0808
		x"00",x"FE",x"01",x"04",x"01",x"FE",x"04",x"04", -- 0x0810
		x"00",x"FE",x"00",x"04",x"04",x"00",x"FE",x"01", -- 0x0818
		x"04",x"FF",x"FE",x"01",x"05",x"00",x"FE",x"05", -- 0x0820
		x"05",x"FF",x"FE",x"01",x"06",x"FF",x"FE",x"01", -- 0x0828
		x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FE",x"01", -- 0x0830
		x"06",x"FE",x"FE",x"01",x"06",x"FE",x"FF",x"01", -- 0x0838
		x"07",x"FE",x"FE",x"05",x"07",x"FE",x"FF",x"01", -- 0x0840
		x"07",x"FE",x"00",x"01",x"08",x"FE",x"FF",x"05", -- 0x0848
		x"08",x"FE",x"00",x"00",x"08",x"00",x"02",x"00", -- 0x0850
		x"01",x"00",x"02",x"FF",x"01",x"01",x"02",x"00", -- 0x0858
		x"06",x"01",x"02",x"FF",x"01",x"01",x"02",x"FE", -- 0x0860
		x"01",x"02",x"02",x"FF",x"03",x"02",x"02",x"FE", -- 0x0868
		x"01",x"02",x"01",x"FE",x"01",x"02",x"02",x"FE", -- 0x0870
		x"02",x"02",x"01",x"FE",x"01",x"03",x"02",x"FE", -- 0x0878
		x"04",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x0880
		x"02",x"03",x"01",x"FE",x"02",x"04",x"00",x"FE", -- 0x0888
		x"01",x"04",x"01",x"FE",x"05",x"04",x"00",x"FE", -- 0x0890
		x"00",x"05",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x0898
		x"FE",x"02",x"04",x"00",x"FE",x"02",x"05",x"FF", -- 0x08A0
		x"FE",x"01",x"05",x"00",x"FE",x"04",x"05",x"FF", -- 0x08A8
		x"FE",x"01",x"05",x"FE",x"FE",x"02",x"06",x"FF", -- 0x08B0
		x"FE",x"01",x"06",x"FE",x"FE",x"01",x"06",x"FF", -- 0x08B8
		x"FE",x"03",x"06",x"FE",x"FE",x"01",x"06",x"FE", -- 0x08C0
		x"FF",x"01",x"07",x"FE",x"FE",x"06",x"07",x"FE", -- 0x08C8
		x"FF",x"01",x"07",x"FE",x"00",x"01",x"08",x"FE", -- 0x08D0
		x"FF",x"08",x"08",x"FE",x"00",x"00",x"0A",x"00", -- 0x08D8
		x"02",x"00",x"01",x"00",x"02",x"FF",x"01",x"01", -- 0x08E0
		x"02",x"00",x"02",x"01",x"02",x"FF",x"01",x"01", -- 0x08E8
		x"02",x"00",x"03",x"01",x"02",x"FF",x"01",x"01", -- 0x08F0
		x"02",x"FE",x"01",x"01",x"02",x"FF",x"01",x"01", -- 0x08F8
		x"02",x"FE",x"01",x"02",x"02",x"FF",x"01",x"02", -- 0x0900
		x"01",x"FE",x"03",x"02",x"02",x"FE",x"02",x"02", -- 0x0908
		x"01",x"FE",x"01",x"02",x"02",x"FE",x"01",x"03", -- 0x0910
		x"02",x"FE",x"01",x"03",x"01",x"FE",x"01",x"03", -- 0x0918
		x"00",x"FE",x"01",x"03",x"02",x"FE",x"01",x"03", -- 0x0920
		x"00",x"FE",x"01",x"03",x"01",x"FE",x"01",x"03", -- 0x0928
		x"00",x"FE",x"01",x"03",x"01",x"FE",x"01",x"03", -- 0x0930
		x"00",x"FE",x"01",x"04",x"01",x"FE",x"02",x"04", -- 0x0938
		x"00",x"FE",x"01",x"04",x"01",x"FE",x"06",x"04", -- 0x0940
		x"00",x"FE",x"01",x"04",x"00",x"FF",x"02",x"04", -- 0x0948
		x"00",x"FE",x"00",x"02",x"04",x"00",x"FE",x"01", -- 0x0950
		x"04",x"00",x"FF",x"06",x"04",x"00",x"FE",x"01", -- 0x0958
		x"04",x"FF",x"FE",x"02",x"04",x"00",x"FE",x"01", -- 0x0960
		x"04",x"FF",x"FE",x"01",x"05",x"00",x"FE",x"01", -- 0x0968
		x"05",x"FF",x"FE",x"01",x"05",x"00",x"FE",x"01", -- 0x0970
		x"05",x"FF",x"FE",x"01",x"05",x"00",x"FE",x"01", -- 0x0978
		x"05",x"FE",x"FE",x"01",x"05",x"00",x"FE",x"01", -- 0x0980
		x"05",x"FF",x"FE",x"01",x"05",x"FE",x"FE",x"01", -- 0x0988
		x"06",x"FE",x"FE",x"02",x"06",x"FF",x"FE",x"03", -- 0x0990
		x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FE",x"01", -- 0x0998
		x"06",x"FE",x"FF",x"01",x"07",x"FE",x"FE",x"01", -- 0x09A0
		x"07",x"FE",x"FF",x"01",x"07",x"FE",x"FE",x"03", -- 0x09A8
		x"07",x"FE",x"FF",x"01",x"07",x"FE",x"00",x"02", -- 0x09B0
		x"07",x"FE",x"FF",x"01",x"07",x"FE",x"00",x"01", -- 0x09B8
		x"08",x"FE",x"FF",x"0A",x"08",x"FE",x"00",x"00", -- 0x09C0
		x"0B",x"00",x"02",x"00",x"01",x"00",x"02",x"FF", -- 0x09C8
		x"01",x"01",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x09D0
		x"01",x"01",x"02",x"00",x"04",x"01",x"02",x"FF", -- 0x09D8
		x"01",x"01",x"02",x"FE",x"01",x"01",x"02",x"FF", -- 0x09E0
		x"02",x"01",x"02",x"FE",x"01",x"02",x"02",x"FF", -- 0x09E8
		x"03",x"02",x"02",x"FE",x"02",x"02",x"01",x"FE", -- 0x09F0
		x"01",x"02",x"02",x"FE",x"02",x"02",x"01",x"FE", -- 0x09F8
		x"01",x"03",x"01",x"FE",x"01",x"03",x"02",x"FE", -- 0x0A00
		x"05",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x0A08
		x"01",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x0A10
		x"01",x"03",x"01",x"FE",x"01",x"04",x"00",x"FE", -- 0x0A18
		x"01",x"04",x"01",x"FE",x"01",x"04",x"00",x"FE", -- 0x0A20
		x"01",x"04",x"01",x"FE",x"06",x"04",x"00",x"FE", -- 0x0A28
		x"00",x"06",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x0A30
		x"FE",x"01",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x0A38
		x"FE",x"01",x"04",x"00",x"FE",x"01",x"05",x"FF", -- 0x0A40
		x"FE",x"01",x"05",x"00",x"FE",x"01",x"05",x"FF", -- 0x0A48
		x"FE",x"01",x"05",x"00",x"FE",x"05",x"05",x"FF", -- 0x0A50
		x"FE",x"01",x"05",x"FE",x"FE",x"01",x"05",x"FF", -- 0x0A58
		x"FE",x"02",x"06",x"FF",x"FE",x"01",x"06",x"FE", -- 0x0A60
		x"FE",x"02",x"06",x"FF",x"FE",x"03",x"06",x"FE", -- 0x0A68
		x"FE",x"01",x"06",x"FE",x"FF",x"02",x"07",x"FE", -- 0x0A70
		x"FE",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x0A78
		x"FE",x"04",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x0A80
		x"00",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x0A88
		x"00",x"01",x"08",x"FE",x"FF",x"0B",x"08",x"FE", -- 0x0A90
		x"00",x"00",x"0B",x"00",x"02",x"00",x"01",x"00", -- 0x0A98
		x"02",x"FF",x"01",x"00",x"02",x"00",x"01",x"01", -- 0x0AA0
		x"02",x"FF",x"01",x"01",x"02",x"00",x"07",x"01", -- 0x0AA8
		x"02",x"FF",x"01",x"01",x"02",x"FE",x"01",x"01", -- 0x0AB0
		x"02",x"FF",x"01",x"01",x"02",x"FE",x"06",x"02", -- 0x0AB8
		x"02",x"FE",x"01",x"02",x"01",x"FE",x"01",x"02", -- 0x0AC0
		x"02",x"FE",x"02",x"02",x"01",x"FE",x"01",x"03", -- 0x0AC8
		x"01",x"FE",x"01",x"03",x"02",x"FE",x"03",x"03", -- 0x0AD0
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"02",x"03", -- 0x0AD8
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"02",x"03", -- 0x0AE0
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"01",x"04", -- 0x0AE8
		x"01",x"FE",x"01",x"04",x"00",x"FE",x"01",x"04", -- 0x0AF0
		x"01",x"FE",x"01",x"04",x"00",x"FE",x"01",x"04", -- 0x0AF8
		x"01",x"FE",x"07",x"04",x"00",x"FE",x"00",x"07", -- 0x0B00
		x"04",x"00",x"FE",x"01",x"04",x"FF",x"FE",x"01", -- 0x0B08
		x"04",x"00",x"FE",x"01",x"04",x"FF",x"FE",x"01", -- 0x0B10
		x"04",x"00",x"FE",x"01",x"04",x"FF",x"FE",x"01", -- 0x0B18
		x"05",x"00",x"FE",x"02",x"05",x"FF",x"FE",x"01", -- 0x0B20
		x"05",x"00",x"FE",x"02",x"05",x"FF",x"FE",x"01", -- 0x0B28
		x"05",x"00",x"FE",x"03",x"05",x"FF",x"FE",x"01", -- 0x0B30
		x"05",x"FE",x"FE",x"01",x"05",x"FF",x"FE",x"02", -- 0x0B38
		x"06",x"FF",x"FE",x"01",x"06",x"FE",x"FE",x"01", -- 0x0B40
		x"06",x"FF",x"FE",x"06",x"06",x"FE",x"FE",x"01", -- 0x0B48
		x"07",x"FE",x"FE",x"01",x"07",x"FE",x"FF",x"01", -- 0x0B50
		x"07",x"FE",x"FE",x"07",x"07",x"FE",x"FF",x"01", -- 0x0B58
		x"07",x"FE",x"00",x"01",x"07",x"FE",x"FF",x"01", -- 0x0B60
		x"08",x"FE",x"00",x"01",x"08",x"FE",x"FF",x"0B", -- 0x0B68
		x"08",x"FE",x"00",x"00",x"0D",x"00",x"02",x"00", -- 0x0B70
		x"01",x"00",x"02",x"FF",x"01",x"01",x"00",x"00", -- 0x0B78
		x"01",x"01",x"02",x"FF",x"01",x"01",x"02",x"00", -- 0x0B80
		x"05",x"01",x"02",x"FF",x"01",x"01",x"02",x"FE", -- 0x0B88
		x"03",x"01",x"02",x"FF",x"02",x"01",x"02",x"FE", -- 0x0B90
		x"02",x"02",x"02",x"FF",x"01",x"02",x"01",x"FE", -- 0x0B98
		x"01",x"02",x"02",x"FF",x"01",x"02",x"01",x"FE", -- 0x0BA0
		x"04",x"02",x"02",x"FE",x"03",x"02",x"01",x"FE", -- 0x0BA8
		x"08",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x0BB0
		x"02",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x0BB8
		x"01",x"03",x"01",x"FE",x"01",x"04",x"00",x"FE", -- 0x0BC0
		x"01",x"04",x"01",x"FE",x"02",x"04",x"00",x"FE", -- 0x0BC8
		x"01",x"04",x"01",x"FE",x"03",x"04",x"00",x"FE", -- 0x0BD0
		x"01",x"04",x"00",x"FF",x"04",x"04",x"00",x"FE", -- 0x0BD8
		x"00",x"04",x"04",x"00",x"FE",x"01",x"04",x"00", -- 0x0BE0
		x"FF",x"03",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x0BE8
		x"FE",x"02",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x0BF0
		x"FE",x"01",x"04",x"00",x"FE",x"01",x"05",x"FF", -- 0x0BF8
		x"FE",x"01",x"05",x"00",x"FE",x"02",x"05",x"FF", -- 0x0C00
		x"FE",x"01",x"05",x"00",x"FE",x"08",x"05",x"FF", -- 0x0C08
		x"FE",x"03",x"06",x"FF",x"FE",x"04",x"06",x"FE", -- 0x0C10
		x"FE",x"01",x"06",x"FF",x"FE",x"01",x"06",x"FE", -- 0x0C18
		x"FF",x"01",x"06",x"FF",x"FE",x"02",x"06",x"FE", -- 0x0C20
		x"FF",x"02",x"07",x"FE",x"FE",x"03",x"07",x"FE", -- 0x0C28
		x"FF",x"01",x"07",x"FE",x"FE",x"05",x"07",x"FE", -- 0x0C30
		x"FF",x"01",x"07",x"FE",x"00",x"01",x"07",x"FE", -- 0x0C38
		x"FF",x"01",x"07",x"00",x"00",x"01",x"08",x"FE", -- 0x0C40
		x"FF",x"0D",x"08",x"FE",x"00",x"00",x"0F",x"00", -- 0x0C48
		x"02",x"00",x"01",x"00",x"02",x"FF",x"03",x"01", -- 0x0C50
		x"02",x"FF",x"01",x"01",x"02",x"00",x"07",x"01", -- 0x0C58
		x"02",x"FF",x"01",x"01",x"02",x"FE",x"01",x"01", -- 0x0C60
		x"02",x"FF",x"01",x"01",x"02",x"FE",x"01",x"02", -- 0x0C68
		x"02",x"FF",x"06",x"02",x"02",x"FE",x"01",x"02", -- 0x0C70
		x"01",x"FE",x"01",x"02",x"02",x"FE",x"02",x"02", -- 0x0C78
		x"01",x"FE",x"01",x"02",x"02",x"FE",x"01",x"02", -- 0x0C80
		x"01",x"FE",x"01",x"03",x"02",x"FE",x"07",x"03", -- 0x0C88
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"02",x"03", -- 0x0C90
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"01",x"03", -- 0x0C98
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"01",x"04", -- 0x0CA0
		x"00",x"FE",x"01",x"04",x"01",x"FE",x"02",x"04", -- 0x0CA8
		x"00",x"FE",x"01",x"04",x"01",x"FE",x"04",x"04", -- 0x0CB0
		x"00",x"FE",x"01",x"04",x"00",x"FF",x"01",x"04", -- 0x0CB8
		x"00",x"FE",x"04",x"04",x"00",x"FE",x"00",x"04", -- 0x0CC0
		x"04",x"00",x"FE",x"01",x"04",x"00",x"FE",x"01", -- 0x0CC8
		x"04",x"00",x"FF",x"04",x"04",x"00",x"FE",x"01", -- 0x0CD0
		x"04",x"FF",x"FE",x"02",x"04",x"00",x"FE",x"01", -- 0x0CD8
		x"04",x"FF",x"FE",x"01",x"04",x"00",x"FE",x"01", -- 0x0CE0
		x"05",x"00",x"FE",x"01",x"05",x"FF",x"FE",x"01", -- 0x0CE8
		x"05",x"00",x"FE",x"02",x"05",x"FF",x"FE",x"01", -- 0x0CF0
		x"05",x"00",x"FE",x"07",x"05",x"FF",x"FE",x"01", -- 0x0CF8
		x"05",x"FE",x"FE",x"01",x"06",x"FF",x"FE",x"01", -- 0x0D00
		x"06",x"FE",x"FE",x"02",x"06",x"FF",x"FE",x"01", -- 0x0D08
		x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FE",x"06", -- 0x0D10
		x"06",x"FE",x"FE",x"01",x"06",x"FE",x"FF",x"01", -- 0x0D18
		x"07",x"FE",x"FE",x"01",x"07",x"FE",x"FF",x"01", -- 0x0D20
		x"07",x"FE",x"FE",x"07",x"07",x"FE",x"FF",x"01", -- 0x0D28
		x"07",x"FE",x"00",x"03",x"07",x"FE",x"FF",x"01", -- 0x0D30
		x"08",x"FE",x"FF",x"0F",x"08",x"FE",x"00",x"00", -- 0x0D38
		x"11",x"00",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x0D40
		x"01",x"01",x"02",x"00",x"03",x"01",x"02",x"FF", -- 0x0D48
		x"01",x"01",x"02",x"00",x"05",x"01",x"02",x"FF", -- 0x0D50
		x"01",x"01",x"02",x"FE",x"01",x"01",x"02",x"FF", -- 0x0D58
		x"01",x"01",x"02",x"FE",x"01",x"01",x"02",x"FF", -- 0x0D60
		x"01",x"01",x"02",x"FE",x"08",x"02",x"02",x"FE", -- 0x0D68
		x"02",x"02",x"01",x"FE",x"01",x"02",x"02",x"FE", -- 0x0D70
		x"01",x"02",x"01",x"FE",x"01",x"02",x"02",x"FE", -- 0x0D78
		x"0A",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x0D80
		x"02",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x0D88
		x"01",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x0D90
		x"01",x"04",x"01",x"FE",x"01",x"04",x"00",x"FE", -- 0x0D98
		x"01",x"04",x"01",x"FE",x"05",x"04",x"00",x"FE", -- 0x0DA0
		x"01",x"04",x"00",x"FF",x"06",x"04",x"00",x"FE", -- 0x0DA8
		x"00",x"06",x"04",x"00",x"FE",x"01",x"04",x"00", -- 0x0DB0
		x"FF",x"05",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x0DB8
		x"FE",x"01",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x0DC0
		x"FE",x"01",x"05",x"00",x"FE",x"01",x"05",x"FF", -- 0x0DC8
		x"FE",x"01",x"05",x"00",x"FE",x"02",x"05",x"FF", -- 0x0DD0
		x"FE",x"01",x"05",x"00",x"FE",x"0A",x"05",x"FF", -- 0x0DD8
		x"FE",x"01",x"06",x"FE",x"FE",x"01",x"06",x"FF", -- 0x0DE0
		x"FE",x"01",x"06",x"FE",x"FE",x"02",x"06",x"FF", -- 0x0DE8
		x"FE",x"08",x"06",x"FE",x"FE",x"01",x"07",x"FE", -- 0x0DF0
		x"FE",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x0DF8
		x"FE",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x0E00
		x"FE",x"05",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x0E08
		x"00",x"03",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x0E10
		x"00",x"01",x"07",x"FE",x"FF",x"11",x"08",x"FE", -- 0x0E18
		x"00",x"00",x"12",x"00",x"02",x"00",x"01",x"00", -- 0x0E20
		x"02",x"FF",x"01",x"01",x"02",x"FF",x"02",x"01", -- 0x0E28
		x"02",x"00",x"03",x"01",x"02",x"FF",x"01",x"01", -- 0x0E30
		x"02",x"00",x"07",x"01",x"02",x"FF",x"01",x"01", -- 0x0E38
		x"02",x"FE",x"01",x"01",x"02",x"FF",x"01",x"01", -- 0x0E40
		x"02",x"FE",x"01",x"01",x"02",x"FF",x"01",x"02", -- 0x0E48
		x"02",x"FE",x"06",x"02",x"02",x"FE",x"01",x"02", -- 0x0E50
		x"01",x"FE",x"01",x"02",x"02",x"FE",x"01",x"02", -- 0x0E58
		x"01",x"FE",x"01",x"02",x"02",x"FE",x"04",x"02", -- 0x0E60
		x"01",x"FE",x"01",x"03",x"02",x"FE",x"07",x"03", -- 0x0E68
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"02",x"03", -- 0x0E70
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"02",x"03", -- 0x0E78
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"01",x"03", -- 0x0E80
		x"01",x"FE",x"01",x"03",x"00",x"FE",x"01",x"04", -- 0x0E88
		x"00",x"FE",x"02",x"04",x"01",x"FE",x"06",x"04", -- 0x0E90
		x"00",x"FE",x"01",x"04",x"00",x"FF",x"06",x"04", -- 0x0E98
		x"00",x"FE",x"00",x"06",x"04",x"00",x"FE",x"01", -- 0x0EA0
		x"04",x"00",x"FF",x"06",x"04",x"00",x"FE",x"02", -- 0x0EA8
		x"04",x"FF",x"FE",x"01",x"04",x"00",x"FE",x"01", -- 0x0EB0
		x"05",x"00",x"FE",x"01",x"05",x"FF",x"FE",x"01", -- 0x0EB8
		x"05",x"00",x"FE",x"02",x"05",x"FF",x"FE",x"01", -- 0x0EC0
		x"05",x"00",x"FE",x"02",x"05",x"FF",x"FE",x"01", -- 0x0EC8
		x"05",x"00",x"FE",x"07",x"05",x"FF",x"FE",x"01", -- 0x0ED0
		x"05",x"FE",x"FE",x"04",x"06",x"FF",x"FE",x"01", -- 0x0ED8
		x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FE",x"01", -- 0x0EE0
		x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FE",x"06", -- 0x0EE8
		x"06",x"FE",x"FE",x"01",x"06",x"FE",x"FE",x"01", -- 0x0EF0
		x"07",x"FE",x"FF",x"01",x"07",x"FE",x"FE",x"01", -- 0x0EF8
		x"07",x"FE",x"FF",x"01",x"07",x"FE",x"FE",x"07", -- 0x0F00
		x"07",x"FE",x"FF",x"01",x"07",x"FE",x"00",x"03", -- 0x0F08
		x"07",x"FE",x"FF",x"02",x"07",x"FE",x"00",x"01", -- 0x0F10
		x"07",x"FE",x"FF",x"01",x"08",x"FE",x"FF",x"12", -- 0x0F18
		x"08",x"FE",x"00",x"00",x"1B",x"00",x"02",x"00", -- 0x0F20
		x"05",x"01",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x0F28
		x"01",x"01",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x0F30
		x"01",x"01",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x0F38
		x"01",x"01",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x0F40
		x"01",x"01",x"02",x"00",x"05",x"01",x"02",x"FF", -- 0x0F48
		x"01",x"01",x"02",x"00",x"04",x"01",x"02",x"FF", -- 0x0F50
		x"01",x"01",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x0F58
		x"01",x"01",x"02",x"FE",x"01",x"01",x"02",x"FF", -- 0x0F60
		x"01",x"01",x"02",x"FE",x"01",x"01",x"02",x"FF", -- 0x0F68
		x"02",x"02",x"02",x"FF",x"01",x"02",x"02",x"FE", -- 0x0F70
		x"01",x"02",x"02",x"FF",x"04",x"02",x"02",x"FE", -- 0x0F78
		x"01",x"02",x"01",x"FE",x"03",x"02",x"02",x"FE", -- 0x0F80
		x"02",x"02",x"01",x"FE",x"01",x"02",x"02",x"FE", -- 0x0F88
		x"04",x"02",x"01",x"FE",x"01",x"02",x"02",x"FE", -- 0x0F90
		x"04",x"02",x"01",x"FE",x"04",x"03",x"01",x"FE", -- 0x0F98
		x"01",x"03",x"00",x"FE",x"04",x"03",x"01",x"FE", -- 0x0FA0
		x"01",x"03",x"00",x"FE",x"02",x"03",x"01",x"FE", -- 0x0FA8
		x"01",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x0FB0
		x"01",x"03",x"00",x"FE",x"02",x"03",x"01",x"FE", -- 0x0FB8
		x"01",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x0FC0
		x"01",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x0FC8
		x"01",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x0FD0
		x"01",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x0FD8
		x"02",x"03",x"00",x"FE",x"01",x"04",x"00",x"FE", -- 0x0FE0
		x"01",x"04",x"01",x"FE",x"06",x"04",x"00",x"FE", -- 0x0FE8
		x"01",x"04",x"01",x"FE",x"07",x"04",x"00",x"FE", -- 0x0FF0
		x"01",x"04",x"00",x"FF",x"08",x"04",x"00",x"FE", -- 0x0FF8
		x"00",x"08",x"04",x"00",x"FE",x"01",x"04",x"00", -- 0x1000
		x"FF",x"07",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x1008
		x"FE",x"06",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x1010
		x"FE",x"01",x"04",x"00",x"FE",x"02",x"05",x"00", -- 0x1018
		x"FE",x"01",x"05",x"FF",x"FE",x"01",x"05",x"00", -- 0x1020
		x"FE",x"01",x"05",x"FF",x"FE",x"01",x"05",x"00", -- 0x1028
		x"FE",x"01",x"05",x"FF",x"FE",x"01",x"05",x"00", -- 0x1030
		x"FE",x"01",x"05",x"FF",x"FE",x"01",x"05",x"00", -- 0x1038
		x"FE",x"02",x"05",x"FF",x"FE",x"01",x"05",x"00", -- 0x1040
		x"FE",x"01",x"05",x"FF",x"FE",x"01",x"05",x"00", -- 0x1048
		x"FE",x"02",x"05",x"FF",x"FE",x"01",x"05",x"00", -- 0x1050
		x"FE",x"04",x"05",x"FF",x"FE",x"01",x"05",x"00", -- 0x1058
		x"FE",x"04",x"05",x"FF",x"FE",x"04",x"06",x"FF", -- 0x1060
		x"FE",x"01",x"06",x"FE",x"FE",x"04",x"06",x"FF", -- 0x1068
		x"FE",x"01",x"06",x"FE",x"FE",x"02",x"06",x"FF", -- 0x1070
		x"FE",x"03",x"06",x"FE",x"FE",x"01",x"06",x"FF", -- 0x1078
		x"FE",x"04",x"06",x"FE",x"FE",x"01",x"06",x"FE", -- 0x1080
		x"FF",x"01",x"06",x"FE",x"FE",x"02",x"06",x"FE", -- 0x1088
		x"FF",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x1090
		x"FE",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x1098
		x"FE",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x10A0
		x"00",x"04",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x10A8
		x"00",x"05",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x10B0
		x"00",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x10B8
		x"00",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x10C0
		x"00",x"01",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x10C8
		x"00",x"01",x"07",x"FE",x"FF",x"05",x"07",x"FE", -- 0x10D0
		x"00",x"1B",x"08",x"FE",x"00",x"00",x"01",x"01", -- 0x10D8
		x"01",x"00",x"02",x"01",x"01",x"00",x"02",x"01", -- 0x10E0
		x"01",x"00",x"02",x"01",x"01",x"00",x"02",x"01", -- 0x10E8
		x"01",x"00",x"02",x"01",x"01",x"00",x"02",x"01", -- 0x10F0
		x"01",x"00",x"02",x"01",x"01",x"00",x"02",x"01", -- 0x10F8
		x"01",x"00",x"02",x"01",x"01",x"00",x"02",x"01", -- 0x1100
		x"08",x"01",x"01",x"01",x"01",x"02",x"01",x"01", -- 0x1108
		x"01",x"02",x"01",x"01",x"01",x"02",x"01",x"01", -- 0x1110
		x"01",x"02",x"01",x"01",x"01",x"02",x"01",x"01", -- 0x1118
		x"01",x"02",x"01",x"01",x"02",x"02",x"01",x"01", -- 0x1120
		x"02",x"02",x"01",x"01",x"02",x"02",x"01",x"01", -- 0x1128
		x"02",x"02",x"01",x"01",x"03",x"02",x"01",x"01", -- 0x1130
		x"03",x"02",x"01",x"01",x"03",x"02",x"01",x"01", -- 0x1138
		x"03",x"02",x"24",x"02",x"00",x"02",x"0C",x"00", -- 0x1140
		x"02",x"01",x"0D",x"01",x"02",x"01",x"0D",x"00", -- 0x1148
		x"02",x"01",x"0D",x"01",x"02",x"01",x"0D",x"00", -- 0x1150
		x"02",x"01",x"0D",x"01",x"02",x"01",x"0D",x"00", -- 0x1158
		x"02",x"06",x"0D",x"01",x"02",x"04",x"0E",x"02", -- 0x1160
		x"02",x"01",x"0E",x"02",x"01",x"01",x"0F",x"02", -- 0x1168
		x"02",x"05",x"0F",x"02",x"01",x"01",x"00",x"02", -- 0x1170
		x"00",x"01",x"00",x"02",x"01",x"01",x"00",x"02", -- 0x1178
		x"00",x"01",x"00",x"02",x"01",x"01",x"00",x"02", -- 0x1180
		x"00",x"01",x"00",x"02",x"01",x"00",x"03",x"00", -- 0x1188
		x"02",x"00",x"01",x"01",x"02",x"FF",x"01",x"01", -- 0x1190
		x"02",x"00",x"01",x"01",x"02",x"FF",x"01",x"01", -- 0x1198
		x"02",x"00",x"01",x"01",x"02",x"FF",x"01",x"01", -- 0x11A0
		x"02",x"00",x"02",x"01",x"02",x"FF",x"01",x"01", -- 0x11A8
		x"02",x"FF",x"01",x"01",x"02",x"00",x"02",x"01", -- 0x11B0
		x"02",x"FF",x"01",x"02",x"02",x"FE",x"01",x"02", -- 0x11B8
		x"02",x"FF",x"08",x"02",x"02",x"FE",x"03",x"02", -- 0x11C0
		x"01",x"FE",x"01",x"02",x"02",x"FE",x"02",x"02", -- 0x11C8
		x"01",x"FE",x"06",x"03",x"01",x"FE",x"01",x"03", -- 0x11D0
		x"00",x"FE",x"01",x"03",x"01",x"FE",x"01",x"03", -- 0x11D8
		x"00",x"FE",x"01",x"03",x"01",x"FE",x"01",x"03", -- 0x11E0
		x"00",x"FE",x"01",x"03",x"01",x"FE",x"01",x"04", -- 0x11E8
		x"00",x"FE",x"01",x"04",x"01",x"FE",x"02",x"04", -- 0x11F0
		x"00",x"FE",x"01",x"04",x"01",x"FE",x"07",x"04", -- 0x11F8
		x"00",x"FE",x"00",x"13",x"92",x"1B",x"92",x"23", -- 0x1200
		x"92",x"2B",x"92",x"33",x"92",x"3B",x"92",x"43", -- 0x1208
		x"92",x"4B",x"92",x"53",x"92",x"94",x"92",x"D5", -- 0x1210
		x"92",x"16",x"93",x"57",x"93",x"B0",x"93",x"09", -- 0x1218
		x"94",x"62",x"94",x"BB",x"94",x"0C",x"95",x"5D", -- 0x1220
		x"95",x"AE",x"95",x"FF",x"95",x"5C",x"96",x"B9", -- 0x1228
		x"96",x"16",x"97",x"73",x"97",x"D4",x"97",x"35", -- 0x1230
		x"98",x"96",x"98",x"F7",x"98",x"68",x"99",x"D9", -- 0x1238
		x"99",x"4A",x"9A",x"BB",x"9A",x"2C",x"9B",x"9D", -- 0x1240
		x"9B",x"0E",x"9C",x"7F",x"9C",x"08",x"9D",x"91", -- 0x1248
		x"9D",x"1A",x"9E",x"07",x"00",x"03",x"00",x"04", -- 0x1250
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x1258
		x"01",x"03",x"FF",x"02",x"01",x"02",x"FE",x"04", -- 0x1260
		x"02",x"02",x"FE",x"02",x"02",x"01",x"FE",x"01", -- 0x1268
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FE",x"01", -- 0x1270
		x"03",x"02",x"FE",x"06",x"03",x"01",x"FD",x"01", -- 0x1278
		x"04",x"00",x"FD",x"01",x"04",x"01",x"FD",x"02", -- 0x1280
		x"04",x"00",x"FD",x"01",x"04",x"00",x"FE",x"01", -- 0x1288
		x"04",x"00",x"FD",x"00",x"01",x"04",x"00",x"FD", -- 0x1290
		x"01",x"04",x"00",x"FE",x"02",x"04",x"00",x"FD", -- 0x1298
		x"01",x"04",x"FF",x"FD",x"01",x"04",x"00",x"FD", -- 0x12A0
		x"06",x"05",x"FF",x"FD",x"01",x"05",x"FE",x"FE", -- 0x12A8
		x"01",x"06",x"FF",x"FE",x"01",x"06",x"FE",x"FE", -- 0x12B0
		x"02",x"06",x"FF",x"FE",x"04",x"06",x"FE",x"FE", -- 0x12B8
		x"02",x"07",x"FE",x"FE",x"01",x"07",x"FD",x"FF", -- 0x12C0
		x"01",x"07",x"FE",x"FE",x"04",x"07",x"FD",x"FF", -- 0x12C8
		x"07",x"08",x"FD",x"00",x"00",x"07",x"08",x"FD", -- 0x12D0
		x"00",x"04",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x12D8
		x"02",x"01",x"09",x"FD",x"01",x"02",x"09",x"FE", -- 0x12E0
		x"02",x"04",x"0A",x"FE",x"02",x"02",x"0A",x"FF", -- 0x12E8
		x"02",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x12F0
		x"02",x"01",x"0B",x"FE",x"02",x"06",x"0B",x"FF", -- 0x12F8
		x"03",x"01",x"0C",x"00",x"03",x"01",x"0C",x"FF", -- 0x1300
		x"03",x"02",x"0C",x"00",x"03",x"01",x"0C",x"00", -- 0x1308
		x"02",x"01",x"0C",x"00",x"03",x"00",x"01",x"0C", -- 0x1310
		x"00",x"03",x"01",x"0C",x"00",x"02",x"02",x"0C", -- 0x1318
		x"00",x"03",x"01",x"0C",x"01",x"03",x"01",x"0C", -- 0x1320
		x"00",x"03",x"06",x"0D",x"01",x"03",x"01",x"0D", -- 0x1328
		x"02",x"02",x"01",x"0E",x"01",x"02",x"01",x"0E", -- 0x1330
		x"02",x"02",x"02",x"0E",x"01",x"02",x"04",x"0E", -- 0x1338
		x"02",x"02",x"02",x"0F",x"02",x"02",x"01",x"0F", -- 0x1340
		x"03",x"01",x"01",x"0F",x"02",x"02",x"04",x"0F", -- 0x1348
		x"03",x"01",x"07",x"00",x"03",x"00",x"00",x"08", -- 0x1350
		x"00",x"03",x"00",x"03",x"01",x"03",x"FF",x"01", -- 0x1358
		x"01",x"02",x"FE",x"01",x"01",x"03",x"FF",x"02", -- 0x1360
		x"01",x"02",x"FE",x"01",x"01",x"03",x"FF",x"04", -- 0x1368
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FE",x"01", -- 0x1370
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FE",x"01", -- 0x1378
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FD",x"01", -- 0x1380
		x"03",x"02",x"FE",x"01",x"03",x"01",x"FD",x"01", -- 0x1388
		x"03",x"02",x"FE",x"05",x"03",x"01",x"FD",x"01", -- 0x1390
		x"04",x"01",x"FD",x"01",x"04",x"00",x"FD",x"01", -- 0x1398
		x"04",x"01",x"FD",x"02",x"04",x"00",x"FD",x"01", -- 0x13A0
		x"04",x"00",x"FE",x"01",x"04",x"00",x"FD",x"00", -- 0x13A8
		x"01",x"04",x"00",x"FD",x"01",x"04",x"00",x"FE", -- 0x13B0
		x"02",x"04",x"00",x"FD",x"01",x"04",x"FF",x"FD", -- 0x13B8
		x"01",x"04",x"00",x"FD",x"01",x"04",x"FF",x"FD", -- 0x13C0
		x"05",x"05",x"FF",x"FD",x"01",x"05",x"FE",x"FE", -- 0x13C8
		x"01",x"05",x"FF",x"FD",x"01",x"05",x"FE",x"FE", -- 0x13D0
		x"01",x"06",x"FF",x"FD",x"01",x"06",x"FE",x"FE", -- 0x13D8
		x"01",x"06",x"FF",x"FE",x"01",x"06",x"FE",x"FE", -- 0x13E0
		x"01",x"06",x"FF",x"FE",x"04",x"06",x"FE",x"FE", -- 0x13E8
		x"01",x"07",x"FD",x"FF",x"02",x"07",x"FE",x"FE", -- 0x13F0
		x"01",x"07",x"FD",x"FF",x"01",x"07",x"FE",x"FE", -- 0x13F8
		x"03",x"07",x"FD",x"FF",x"08",x"08",x"FD",x"00", -- 0x1400
		x"00",x"08",x"08",x"FD",x"00",x"03",x"09",x"FD", -- 0x1408
		x"01",x"01",x"09",x"FE",x"02",x"01",x"09",x"FD", -- 0x1410
		x"01",x"02",x"09",x"FE",x"02",x"01",x"09",x"FD", -- 0x1418
		x"01",x"04",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1420
		x"02",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1428
		x"02",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1430
		x"03",x"01",x"0B",x"FE",x"02",x"01",x"0B",x"FF", -- 0x1438
		x"03",x"01",x"0B",x"FE",x"02",x"05",x"0B",x"FF", -- 0x1440
		x"03",x"01",x"0C",x"FF",x"03",x"01",x"0C",x"00", -- 0x1448
		x"03",x"01",x"0C",x"FF",x"03",x"02",x"0C",x"00", -- 0x1450
		x"03",x"01",x"0C",x"00",x"02",x"01",x"0C",x"00", -- 0x1458
		x"03",x"00",x"01",x"0C",x"00",x"03",x"01",x"0C", -- 0x1460
		x"00",x"02",x"02",x"0C",x"00",x"03",x"01",x"0C", -- 0x1468
		x"01",x"03",x"01",x"0C",x"00",x"03",x"01",x"0C", -- 0x1470
		x"01",x"03",x"05",x"0D",x"01",x"03",x"01",x"0D", -- 0x1478
		x"02",x"02",x"01",x"0D",x"01",x"03",x"01",x"0D", -- 0x1480
		x"02",x"02",x"01",x"0E",x"01",x"03",x"01",x"0E", -- 0x1488
		x"02",x"02",x"01",x"0E",x"01",x"02",x"01",x"0E", -- 0x1490
		x"02",x"02",x"01",x"0E",x"01",x"02",x"04",x"0E", -- 0x1498
		x"02",x"02",x"01",x"0F",x"03",x"01",x"02",x"0F", -- 0x14A0
		x"02",x"02",x"01",x"0F",x"03",x"01",x"01",x"0F", -- 0x14A8
		x"02",x"02",x"03",x"0F",x"03",x"01",x"08",x"00", -- 0x14B0
		x"03",x"00",x"00",x"06",x"00",x"03",x"00",x"01", -- 0x14B8
		x"00",x"03",x"FF",x"02",x"00",x"03",x"00",x"03", -- 0x14C0
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x14C8
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FF",x"02", -- 0x14D0
		x"01",x"02",x"FE",x"01",x"01",x"03",x"FF",x"06", -- 0x14D8
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FD",x"01", -- 0x14E0
		x"02",x"02",x"FE",x"02",x"02",x"01",x"FE",x"01", -- 0x14E8
		x"03",x"02",x"FE",x"02",x"03",x"01",x"FD",x"01", -- 0x14F0
		x"03",x"02",x"FE",x"04",x"03",x"01",x"FD",x"01", -- 0x14F8
		x"03",x"00",x"FD",x"03",x"04",x"01",x"FD",x"04", -- 0x1500
		x"04",x"00",x"FD",x"00",x"04",x"04",x"00",x"FD", -- 0x1508
		x"03",x"04",x"FF",x"FD",x"01",x"05",x"00",x"FD", -- 0x1510
		x"04",x"05",x"FF",x"FD",x"01",x"05",x"FE",x"FE", -- 0x1518
		x"02",x"05",x"FF",x"FD",x"01",x"05",x"FE",x"FE", -- 0x1520
		x"02",x"06",x"FF",x"FE",x"01",x"06",x"FE",x"FE", -- 0x1528
		x"01",x"06",x"FF",x"FD",x"06",x"06",x"FE",x"FE", -- 0x1530
		x"01",x"07",x"FD",x"FF",x"02",x"07",x"FE",x"FE", -- 0x1538
		x"01",x"07",x"FE",x"FF",x"01",x"07",x"FD",x"FF", -- 0x1540
		x"01",x"07",x"FE",x"FE",x"03",x"07",x"FD",x"FF", -- 0x1548
		x"02",x"08",x"FD",x"00",x"01",x"08",x"FD",x"FF", -- 0x1550
		x"06",x"08",x"FD",x"00",x"00",x"06",x"08",x"FD", -- 0x1558
		x"00",x"01",x"08",x"FD",x"01",x"02",x"08",x"FD", -- 0x1560
		x"00",x"03",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x1568
		x"02",x"01",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x1570
		x"01",x"02",x"09",x"FE",x"02",x"01",x"09",x"FD", -- 0x1578
		x"01",x"06",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1580
		x"03",x"01",x"0A",x"FE",x"02",x"02",x"0A",x"FF", -- 0x1588
		x"02",x"01",x"0B",x"FE",x"02",x"02",x"0B",x"FF", -- 0x1590
		x"03",x"01",x"0B",x"FE",x"02",x"04",x"0B",x"FF", -- 0x1598
		x"03",x"01",x"0B",x"00",x"03",x"03",x"0C",x"FF", -- 0x15A0
		x"03",x"04",x"0C",x"00",x"03",x"00",x"04",x"0C", -- 0x15A8
		x"00",x"03",x"03",x"0C",x"01",x"03",x"01",x"0D", -- 0x15B0
		x"00",x"03",x"04",x"0D",x"01",x"03",x"01",x"0D", -- 0x15B8
		x"02",x"02",x"02",x"0D",x"01",x"03",x"01",x"0D", -- 0x15C0
		x"02",x"02",x"02",x"0E",x"01",x"02",x"01",x"0E", -- 0x15C8
		x"02",x"02",x"01",x"0E",x"01",x"03",x"06",x"0E", -- 0x15D0
		x"02",x"02",x"01",x"0F",x"03",x"01",x"02",x"0F", -- 0x15D8
		x"02",x"02",x"01",x"0F",x"02",x"01",x"01",x"0F", -- 0x15E0
		x"03",x"01",x"01",x"0F",x"02",x"02",x"03",x"0F", -- 0x15E8
		x"03",x"01",x"02",x"00",x"03",x"00",x"01",x"00", -- 0x15F0
		x"03",x"01",x"06",x"00",x"03",x"00",x"00",x"08", -- 0x15F8
		x"00",x"03",x"00",x"02",x"00",x"03",x"FF",x"03", -- 0x1600
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x1608
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x1610
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x1618
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"08", -- 0x1620
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FD",x"01", -- 0x1628
		x"02",x"02",x"FE",x"01",x"03",x"01",x"FD",x"01", -- 0x1630
		x"03",x"02",x"FE",x"04",x"03",x"01",x"FD",x"01", -- 0x1638
		x"03",x"02",x"FE",x"01",x"03",x"00",x"FD",x"02", -- 0x1640
		x"03",x"01",x"FD",x"01",x"04",x"01",x"FD",x"01", -- 0x1648
		x"04",x"00",x"FD",x"01",x"04",x"01",x"FD",x"05", -- 0x1650
		x"04",x"00",x"FD",x"00",x"05",x"04",x"00",x"FD", -- 0x1658
		x"01",x"04",x"FF",x"FD",x"01",x"04",x"00",x"FD", -- 0x1660
		x"01",x"04",x"FF",x"FD",x"02",x"05",x"FF",x"FD", -- 0x1668
		x"01",x"05",x"00",x"FD",x"01",x"05",x"FE",x"FE", -- 0x1670
		x"04",x"05",x"FF",x"FD",x"01",x"05",x"FE",x"FE", -- 0x1678
		x"01",x"05",x"FF",x"FD",x"01",x"06",x"FE",x"FE", -- 0x1680
		x"01",x"06",x"FF",x"FD",x"08",x"06",x"FE",x"FE", -- 0x1688
		x"01",x"07",x"FE",x"FE",x"01",x"07",x"FD",x"FF", -- 0x1690
		x"01",x"07",x"FE",x"FE",x"01",x"07",x"FD",x"FF", -- 0x1698
		x"01",x"07",x"FE",x"FE",x"01",x"07",x"FD",x"FF", -- 0x16A0
		x"01",x"07",x"FE",x"FE",x"03",x"07",x"FD",x"FF", -- 0x16A8
		x"02",x"08",x"FD",x"FF",x"08",x"08",x"FD",x"00", -- 0x16B0
		x"00",x"08",x"08",x"FD",x"00",x"02",x"08",x"FD", -- 0x16B8
		x"01",x"03",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x16C0
		x"02",x"01",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x16C8
		x"02",x"01",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x16D0
		x"02",x"01",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x16D8
		x"02",x"08",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x16E0
		x"03",x"01",x"0A",x"FE",x"02",x"01",x"0B",x"FF", -- 0x16E8
		x"03",x"01",x"0B",x"FE",x"02",x"04",x"0B",x"FF", -- 0x16F0
		x"03",x"01",x"0B",x"FE",x"02",x"01",x"0B",x"00", -- 0x16F8
		x"03",x"02",x"0B",x"FF",x"03",x"01",x"0C",x"FF", -- 0x1700
		x"03",x"01",x"0C",x"00",x"03",x"01",x"0C",x"FF", -- 0x1708
		x"03",x"05",x"0C",x"00",x"03",x"00",x"05",x"0C", -- 0x1710
		x"00",x"03",x"01",x"0C",x"01",x"03",x"01",x"0C", -- 0x1718
		x"00",x"03",x"01",x"0C",x"01",x"03",x"02",x"0D", -- 0x1720
		x"01",x"03",x"01",x"0D",x"00",x"03",x"01",x"0D", -- 0x1728
		x"02",x"02",x"04",x"0D",x"01",x"03",x"01",x"0D", -- 0x1730
		x"02",x"02",x"01",x"0D",x"01",x"03",x"01",x"0E", -- 0x1738
		x"02",x"02",x"01",x"0E",x"01",x"03",x"08",x"0E", -- 0x1740
		x"02",x"02",x"01",x"0F",x"02",x"02",x"01",x"0F", -- 0x1748
		x"03",x"01",x"01",x"0F",x"02",x"02",x"01",x"0F", -- 0x1750
		x"03",x"01",x"01",x"0F",x"02",x"02",x"01",x"0F", -- 0x1758
		x"03",x"01",x"01",x"0F",x"02",x"02",x"03",x"0F", -- 0x1760
		x"03",x"01",x"02",x"00",x"03",x"01",x"08",x"00", -- 0x1768
		x"03",x"00",x"00",x"09",x"00",x"03",x"00",x"01", -- 0x1770
		x"00",x"03",x"FF",x"06",x"01",x"03",x"FF",x"01", -- 0x1778
		x"01",x"02",x"FE",x"01",x"01",x"03",x"FF",x"01", -- 0x1780
		x"01",x"02",x"FE",x"01",x"01",x"03",x"FF",x"02", -- 0x1788
		x"01",x"02",x"FE",x"07",x"02",x"02",x"FE",x"02", -- 0x1790
		x"02",x"01",x"FE",x"01",x"02",x"02",x"FE",x"01", -- 0x1798
		x"02",x"01",x"FE",x"01",x"02",x"02",x"FE",x"01", -- 0x17A0
		x"03",x"01",x"FD",x"01",x"03",x"02",x"FE",x"02", -- 0x17A8
		x"03",x"01",x"FD",x"01",x"03",x"01",x"FE",x"01", -- 0x17B0
		x"03",x"01",x"FD",x"01",x"03",x"01",x"FE",x"03", -- 0x17B8
		x"03",x"01",x"FD",x"01",x"04",x"01",x"FD",x"01", -- 0x17C0
		x"04",x"00",x"FD",x"01",x"04",x"01",x"FD",x"06", -- 0x17C8
		x"04",x"00",x"FD",x"00",x"06",x"04",x"00",x"FD", -- 0x17D0
		x"01",x"04",x"FF",x"FD",x"01",x"04",x"00",x"FD", -- 0x17D8
		x"01",x"04",x"FF",x"FD",x"03",x"05",x"FF",x"FD", -- 0x17E0
		x"01",x"05",x"FF",x"FE",x"01",x"05",x"FF",x"FD", -- 0x17E8
		x"01",x"05",x"FF",x"FE",x"02",x"05",x"FF",x"FD", -- 0x17F0
		x"01",x"05",x"FE",x"FE",x"01",x"05",x"FF",x"FD", -- 0x17F8
		x"01",x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FE", -- 0x1800
		x"01",x"06",x"FE",x"FE",x"02",x"06",x"FF",x"FE", -- 0x1808
		x"07",x"06",x"FE",x"FE",x"02",x"07",x"FE",x"FE", -- 0x1810
		x"01",x"07",x"FD",x"FF",x"01",x"07",x"FE",x"FE", -- 0x1818
		x"01",x"07",x"FD",x"FF",x"01",x"07",x"FE",x"FE", -- 0x1820
		x"06",x"07",x"FD",x"FF",x"01",x"08",x"FD",x"FF", -- 0x1828
		x"09",x"08",x"FD",x"00",x"00",x"09",x"08",x"FD", -- 0x1830
		x"00",x"01",x"08",x"FD",x"01",x"06",x"09",x"FD", -- 0x1838
		x"01",x"01",x"09",x"FE",x"02",x"01",x"09",x"FD", -- 0x1840
		x"01",x"01",x"09",x"FE",x"02",x"01",x"09",x"FD", -- 0x1848
		x"01",x"02",x"09",x"FE",x"02",x"07",x"0A",x"FE", -- 0x1850
		x"02",x"02",x"0A",x"FF",x"02",x"01",x"0A",x"FE", -- 0x1858
		x"02",x"01",x"0A",x"FF",x"02",x"01",x"0A",x"FE", -- 0x1860
		x"02",x"01",x"0B",x"FF",x"03",x"01",x"0B",x"FE", -- 0x1868
		x"02",x"02",x"0B",x"FF",x"03",x"01",x"0B",x"FF", -- 0x1870
		x"02",x"01",x"0B",x"FF",x"03",x"01",x"0B",x"FF", -- 0x1878
		x"02",x"03",x"0B",x"FF",x"03",x"01",x"0C",x"FF", -- 0x1880
		x"03",x"01",x"0C",x"00",x"03",x"01",x"0C",x"FF", -- 0x1888
		x"03",x"06",x"0C",x"00",x"03",x"00",x"06",x"0C", -- 0x1890
		x"00",x"03",x"01",x"0C",x"01",x"03",x"01",x"0C", -- 0x1898
		x"00",x"03",x"01",x"0C",x"01",x"03",x"03",x"0D", -- 0x18A0
		x"01",x"03",x"01",x"0D",x"01",x"02",x"01",x"0D", -- 0x18A8
		x"01",x"03",x"01",x"0D",x"01",x"02",x"02",x"0D", -- 0x18B0
		x"01",x"03",x"01",x"0D",x"02",x"02",x"01",x"0D", -- 0x18B8
		x"01",x"03",x"01",x"0E",x"02",x"02",x"01",x"0E", -- 0x18C0
		x"01",x"02",x"01",x"0E",x"02",x"02",x"02",x"0E", -- 0x18C8
		x"01",x"02",x"07",x"0E",x"02",x"02",x"02",x"0F", -- 0x18D0
		x"02",x"02",x"01",x"0F",x"03",x"01",x"01",x"0F", -- 0x18D8
		x"02",x"02",x"01",x"0F",x"03",x"01",x"01",x"0F", -- 0x18E0
		x"02",x"02",x"06",x"0F",x"03",x"01",x"01",x"00", -- 0x18E8
		x"03",x"01",x"09",x"00",x"03",x"00",x"00",x"0B", -- 0x18F0
		x"00",x"03",x"00",x"01",x"01",x"03",x"FF",x"01", -- 0x18F8
		x"01",x"03",x"00",x"02",x"01",x"03",x"FF",x"01", -- 0x1900
		x"01",x"02",x"FE",x"02",x"01",x"03",x"FF",x"01", -- 0x1908
		x"01",x"02",x"FE",x"01",x"01",x"03",x"FF",x"03", -- 0x1910
		x"01",x"02",x"FE",x"01",x"01",x"03",x"FF",x"05", -- 0x1918
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FE",x"02", -- 0x1920
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FE",x"01", -- 0x1928
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FD",x"01", -- 0x1930
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FE",x"01", -- 0x1938
		x"03",x"02",x"FE",x"02",x"03",x"01",x"FD",x"01", -- 0x1940
		x"03",x"02",x"FE",x"03",x"03",x"01",x"FD",x"02", -- 0x1948
		x"03",x"01",x"FE",x"02",x"03",x"01",x"FD",x"01", -- 0x1950
		x"04",x"01",x"FD",x"01",x"04",x"00",x"FD",x"01", -- 0x1958
		x"04",x"01",x"FD",x"07",x"04",x"00",x"FD",x"00", -- 0x1960
		x"07",x"04",x"00",x"FD",x"01",x"04",x"FF",x"FD", -- 0x1968
		x"01",x"04",x"00",x"FD",x"01",x"04",x"FF",x"FD", -- 0x1970
		x"02",x"05",x"FF",x"FD",x"02",x"05",x"FF",x"FE", -- 0x1978
		x"03",x"05",x"FF",x"FD",x"01",x"05",x"FE",x"FE", -- 0x1980
		x"02",x"05",x"FF",x"FD",x"01",x"05",x"FE",x"FE", -- 0x1988
		x"01",x"06",x"FF",x"FE",x"01",x"06",x"FE",x"FE", -- 0x1990
		x"01",x"06",x"FF",x"FD",x"01",x"06",x"FE",x"FE", -- 0x1998
		x"01",x"06",x"FF",x"FE",x"02",x"06",x"FE",x"FE", -- 0x19A0
		x"01",x"06",x"FF",x"FE",x"05",x"06",x"FE",x"FE", -- 0x19A8
		x"01",x"07",x"FD",x"FF",x"03",x"07",x"FE",x"FE", -- 0x19B0
		x"01",x"07",x"FD",x"FF",x"01",x"07",x"FE",x"FE", -- 0x19B8
		x"02",x"07",x"FD",x"FF",x"01",x"07",x"FE",x"FE", -- 0x19C0
		x"02",x"07",x"FD",x"FF",x"01",x"07",x"FD",x"00", -- 0x19C8
		x"01",x"07",x"FD",x"FF",x"0B",x"08",x"FD",x"00", -- 0x19D0
		x"00",x"0B",x"08",x"FD",x"00",x"01",x"09",x"FD", -- 0x19D8
		x"01",x"01",x"09",x"FD",x"00",x"02",x"09",x"FD", -- 0x19E0
		x"01",x"01",x"09",x"FE",x"02",x"02",x"09",x"FD", -- 0x19E8
		x"01",x"01",x"09",x"FE",x"02",x"01",x"09",x"FD", -- 0x19F0
		x"01",x"03",x"09",x"FE",x"02",x"01",x"09",x"FD", -- 0x19F8
		x"01",x"05",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1A00
		x"02",x"02",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1A08
		x"02",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1A10
		x"03",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1A18
		x"02",x"01",x"0B",x"FE",x"02",x"02",x"0B",x"FF", -- 0x1A20
		x"03",x"01",x"0B",x"FE",x"02",x"03",x"0B",x"FF", -- 0x1A28
		x"03",x"02",x"0B",x"FF",x"02",x"02",x"0B",x"FF", -- 0x1A30
		x"03",x"01",x"0C",x"FF",x"03",x"01",x"0C",x"00", -- 0x1A38
		x"03",x"01",x"0C",x"FF",x"03",x"07",x"0C",x"00", -- 0x1A40
		x"03",x"00",x"07",x"0C",x"00",x"03",x"01",x"0C", -- 0x1A48
		x"01",x"03",x"01",x"0C",x"00",x"03",x"01",x"0C", -- 0x1A50
		x"01",x"03",x"02",x"0D",x"01",x"03",x"02",x"0D", -- 0x1A58
		x"01",x"02",x"03",x"0D",x"01",x"03",x"01",x"0D", -- 0x1A60
		x"02",x"02",x"02",x"0D",x"01",x"03",x"01",x"0D", -- 0x1A68
		x"02",x"02",x"01",x"0E",x"01",x"02",x"01",x"0E", -- 0x1A70
		x"02",x"02",x"01",x"0E",x"01",x"03",x"01",x"0E", -- 0x1A78
		x"02",x"02",x"01",x"0E",x"01",x"02",x"02",x"0E", -- 0x1A80
		x"02",x"02",x"01",x"0E",x"01",x"02",x"05",x"0E", -- 0x1A88
		x"02",x"02",x"01",x"0F",x"03",x"01",x"03",x"0F", -- 0x1A90
		x"02",x"02",x"01",x"0F",x"03",x"01",x"01",x"0F", -- 0x1A98
		x"02",x"02",x"02",x"0F",x"03",x"01",x"01",x"0F", -- 0x1AA0
		x"02",x"02",x"02",x"0F",x"03",x"01",x"01",x"0F", -- 0x1AA8
		x"03",x"00",x"01",x"0F",x"03",x"01",x"0B",x"00", -- 0x1AB0
		x"03",x"00",x"00",x"0B",x"00",x"03",x"00",x"02", -- 0x1AB8
		x"01",x"03",x"FF",x"01",x"01",x"03",x"00",x"04", -- 0x1AC0
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x1AC8
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x1AD0
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x1AD8
		x"01",x"02",x"FF",x"01",x"01",x"02",x"FE",x"01", -- 0x1AE0
		x"01",x"03",x"FF",x"06",x"02",x"02",x"FE",x"01", -- 0x1AE8
		x"02",x"01",x"FE",x"02",x"02",x"02",x"FE",x"01", -- 0x1AF0
		x"02",x"01",x"FD",x"01",x"02",x"02",x"FE",x"01", -- 0x1AF8
		x"02",x"01",x"FD",x"01",x"03",x"02",x"FE",x"01", -- 0x1B00
		x"03",x"01",x"FD",x"02",x"03",x"02",x"FE",x"01", -- 0x1B08
		x"03",x"01",x"FD",x"07",x"03",x"02",x"FE",x"01", -- 0x1B10
		x"04",x"01",x"FD",x"02",x"04",x"00",x"FD",x"05", -- 0x1B18
		x"04",x"01",x"FD",x"01",x"04",x"00",x"FE",x"02", -- 0x1B20
		x"04",x"00",x"FD",x"00",x"02",x"04",x"00",x"FD", -- 0x1B28
		x"01",x"04",x"00",x"FE",x"05",x"04",x"FF",x"FD", -- 0x1B30
		x"02",x"04",x"00",x"FD",x"01",x"04",x"FF",x"FD", -- 0x1B38
		x"07",x"05",x"FE",x"FE",x"01",x"05",x"FF",x"FD", -- 0x1B40
		x"02",x"05",x"FE",x"FE",x"01",x"05",x"FF",x"FD", -- 0x1B48
		x"01",x"05",x"FE",x"FE",x"01",x"06",x"FF",x"FD", -- 0x1B50
		x"01",x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FD", -- 0x1B58
		x"02",x"06",x"FE",x"FE",x"01",x"06",x"FF",x"FE", -- 0x1B60
		x"06",x"06",x"FE",x"FE",x"01",x"07",x"FD",x"FF", -- 0x1B68
		x"01",x"07",x"FE",x"FE",x"01",x"07",x"FE",x"FF", -- 0x1B70
		x"01",x"07",x"FE",x"FE",x"01",x"07",x"FD",x"FF", -- 0x1B78
		x"01",x"07",x"FE",x"FE",x"01",x"07",x"FD",x"FF", -- 0x1B80
		x"01",x"07",x"FE",x"FE",x"04",x"07",x"FD",x"FF", -- 0x1B88
		x"01",x"07",x"FD",x"00",x"02",x"07",x"FD",x"FF", -- 0x1B90
		x"0B",x"08",x"FD",x"00",x"00",x"0B",x"08",x"FD", -- 0x1B98
		x"00",x"02",x"09",x"FD",x"01",x"01",x"09",x"FD", -- 0x1BA0
		x"00",x"04",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x1BA8
		x"02",x"01",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x1BB0
		x"02",x"01",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x1BB8
		x"02",x"01",x"09",x"FE",x"01",x"01",x"09",x"FE", -- 0x1BC0
		x"02",x"01",x"09",x"FD",x"01",x"06",x"0A",x"FE", -- 0x1BC8
		x"02",x"01",x"0A",x"FF",x"02",x"02",x"0A",x"FE", -- 0x1BD0
		x"02",x"01",x"0A",x"FF",x"03",x"01",x"0A",x"FE", -- 0x1BD8
		x"02",x"01",x"0A",x"FF",x"03",x"01",x"0B",x"FE", -- 0x1BE0
		x"02",x"01",x"0B",x"FF",x"03",x"02",x"0B",x"FE", -- 0x1BE8
		x"02",x"01",x"0B",x"FF",x"03",x"07",x"0B",x"FE", -- 0x1BF0
		x"02",x"01",x"0C",x"FF",x"03",x"02",x"0C",x"00", -- 0x1BF8
		x"03",x"05",x"0C",x"FF",x"03",x"01",x"0C",x"00", -- 0x1C00
		x"02",x"02",x"0C",x"00",x"03",x"00",x"02",x"0C", -- 0x1C08
		x"00",x"03",x"01",x"0C",x"00",x"02",x"05",x"0C", -- 0x1C10
		x"01",x"03",x"02",x"0C",x"00",x"03",x"01",x"0C", -- 0x1C18
		x"01",x"03",x"07",x"0D",x"02",x"02",x"01",x"0D", -- 0x1C20
		x"01",x"03",x"02",x"0D",x"02",x"02",x"01",x"0D", -- 0x1C28
		x"01",x"03",x"01",x"0D",x"02",x"02",x"01",x"0E", -- 0x1C30
		x"01",x"03",x"01",x"0E",x"02",x"02",x"01",x"0E", -- 0x1C38
		x"01",x"03",x"02",x"0E",x"02",x"02",x"01",x"0E", -- 0x1C40
		x"01",x"02",x"06",x"0E",x"02",x"02",x"01",x"0F", -- 0x1C48
		x"03",x"01",x"01",x"0F",x"02",x"02",x"01",x"0F", -- 0x1C50
		x"02",x"01",x"01",x"0F",x"02",x"02",x"01",x"0F", -- 0x1C58
		x"03",x"01",x"01",x"0F",x"02",x"02",x"01",x"0F", -- 0x1C60
		x"03",x"01",x"01",x"0F",x"02",x"02",x"04",x"0F", -- 0x1C68
		x"03",x"01",x"01",x"0F",x"03",x"00",x"02",x"0F", -- 0x1C70
		x"03",x"01",x"0B",x"00",x"03",x"00",x"00",x"12", -- 0x1C78
		x"00",x"03",x"00",x"03",x"01",x"03",x"00",x"02", -- 0x1C80
		x"01",x"03",x"FF",x"01",x"01",x"03",x"00",x"06", -- 0x1C88
		x"01",x"03",x"FF",x"01",x"01",x"02",x"FE",x"04", -- 0x1C90
		x"01",x"03",x"FF",x"03",x"01",x"02",x"FE",x"01", -- 0x1C98
		x"01",x"02",x"FF",x"01",x"02",x"02",x"FF",x"01", -- 0x1CA0
		x"02",x"02",x"FE",x"01",x"02",x"03",x"FF",x"01", -- 0x1CA8
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FE",x"06", -- 0x1CB0
		x"02",x"02",x"FE",x"02",x"02",x"01",x"FE",x"01", -- 0x1CB8
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FD",x"01", -- 0x1CC0
		x"02",x"02",x"FE",x"01",x"02",x"01",x"FD",x"01", -- 0x1CC8
		x"02",x"02",x"FE",x"02",x"02",x"01",x"FE",x"01", -- 0x1CD0
		x"02",x"02",x"FE",x"02",x"02",x"01",x"FD",x"01", -- 0x1CD8
		x"03",x"01",x"FD",x"01",x"03",x"02",x"FE",x"0D", -- 0x1CE0
		x"03",x"01",x"FD",x"01",x"03",x"00",x"FD",x"01", -- 0x1CE8
		x"03",x"01",x"FD",x"01",x"03",x"00",x"FD",x"01", -- 0x1CF0
		x"04",x"01",x"FD",x"04",x"04",x"00",x"FD",x"01", -- 0x1CF8
		x"04",x"01",x"FD",x"0A",x"04",x"00",x"FD",x"00", -- 0x1D00
		x"0A",x"04",x"00",x"FD",x"01",x"04",x"FF",x"FD", -- 0x1D08
		x"04",x"04",x"00",x"FD",x"01",x"04",x"FF",x"FD", -- 0x1D10
		x"01",x"05",x"00",x"FD",x"01",x"05",x"FF",x"FD", -- 0x1D18
		x"01",x"05",x"00",x"FD",x"0D",x"05",x"FF",x"FD", -- 0x1D20
		x"01",x"05",x"FE",x"FE",x"01",x"05",x"FF",x"FD", -- 0x1D28
		x"02",x"06",x"FF",x"FD",x"01",x"06",x"FE",x"FE", -- 0x1D30
		x"02",x"06",x"FF",x"FE",x"01",x"06",x"FE",x"FE", -- 0x1D38
		x"01",x"06",x"FF",x"FD",x"01",x"06",x"FE",x"FE", -- 0x1D40
		x"01",x"06",x"FF",x"FD",x"01",x"06",x"FE",x"FE", -- 0x1D48
		x"02",x"06",x"FF",x"FE",x"06",x"06",x"FE",x"FE", -- 0x1D50
		x"01",x"06",x"FF",x"FE",x"01",x"06",x"FE",x"FE", -- 0x1D58
		x"01",x"06",x"FD",x"FF",x"01",x"06",x"FE",x"FE", -- 0x1D60
		x"01",x"06",x"FE",x"FF",x"01",x"07",x"FE",x"FF", -- 0x1D68
		x"03",x"07",x"FE",x"FE",x"04",x"07",x"FD",x"FF", -- 0x1D70
		x"01",x"07",x"FE",x"FE",x"06",x"07",x"FD",x"FF", -- 0x1D78
		x"01",x"07",x"FD",x"00",x"02",x"07",x"FD",x"FF", -- 0x1D80
		x"03",x"07",x"FD",x"00",x"12",x"08",x"FD",x"00", -- 0x1D88
		x"00",x"12",x"08",x"FD",x"00",x"03",x"09",x"FD", -- 0x1D90
		x"00",x"02",x"09",x"FD",x"01",x"01",x"09",x"FD", -- 0x1D98
		x"00",x"06",x"09",x"FD",x"01",x"01",x"09",x"FE", -- 0x1DA0
		x"02",x"04",x"09",x"FD",x"01",x"03",x"09",x"FE", -- 0x1DA8
		x"02",x"01",x"09",x"FE",x"01",x"01",x"0A",x"FE", -- 0x1DB0
		x"01",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FD", -- 0x1DB8
		x"01",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1DC0
		x"02",x"06",x"0A",x"FE",x"02",x"02",x"0A",x"FF", -- 0x1DC8
		x"02",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1DD0
		x"03",x"01",x"0A",x"FE",x"02",x"01",x"0A",x"FF", -- 0x1DD8
		x"03",x"01",x"0A",x"FE",x"02",x"02",x"0A",x"FF", -- 0x1DE0
		x"02",x"01",x"0A",x"FE",x"02",x"02",x"0A",x"FF", -- 0x1DE8
		x"03",x"01",x"0B",x"FF",x"03",x"01",x"0B",x"FE", -- 0x1DF0
		x"02",x"0D",x"0B",x"FF",x"03",x"01",x"0B",x"00", -- 0x1DF8
		x"03",x"01",x"0B",x"FF",x"03",x"01",x"0B",x"00", -- 0x1E00
		x"03",x"01",x"0C",x"FF",x"03",x"04",x"0C",x"00", -- 0x1E08
		x"03",x"01",x"0C",x"FF",x"03",x"0A",x"0C",x"00", -- 0x1E10
		x"03",x"00",x"0A",x"0C",x"00",x"03",x"01",x"0C", -- 0x1E18
		x"01",x"03",x"04",x"0C",x"00",x"03",x"01",x"0C", -- 0x1E20
		x"01",x"03",x"01",x"0D",x"00",x"03",x"01",x"0D", -- 0x1E28
		x"01",x"03",x"01",x"0D",x"00",x"03",x"0D",x"0D", -- 0x1E30
		x"01",x"03",x"01",x"0D",x"02",x"02",x"01",x"0D", -- 0x1E38
		x"01",x"03",x"02",x"0E",x"01",x"03",x"01",x"0E", -- 0x1E40
		x"02",x"02",x"02",x"0E",x"01",x"02",x"01",x"0E", -- 0x1E48
		x"02",x"02",x"01",x"0E",x"01",x"03",x"01",x"0E", -- 0x1E50
		x"02",x"02",x"01",x"0E",x"01",x"03",x"01",x"0E", -- 0x1E58
		x"02",x"02",x"02",x"0E",x"01",x"02",x"06",x"0E", -- 0x1E60
		x"02",x"02",x"01",x"0E",x"01",x"02",x"01",x"0E", -- 0x1E68
		x"02",x"02",x"01",x"0E",x"03",x"01",x"01",x"0E", -- 0x1E70
		x"02",x"02",x"01",x"0E",x"02",x"01",x"01",x"0F", -- 0x1E78
		x"02",x"01",x"03",x"0F",x"02",x"02",x"04",x"0F", -- 0x1E80
		x"03",x"01",x"01",x"0F",x"02",x"02",x"06",x"0F", -- 0x1E88
		x"03",x"01",x"01",x"0F",x"03",x"00",x"02",x"0F", -- 0x1E90
		x"03",x"01",x"03",x"0F",x"03",x"00",x"12",x"00", -- 0x1E98
		x"03",x"00",x"00",x"00",x"01",x"02",x"02",x"02", -- 0x1EA0
		x"02",x"02",x"02",x"00",x"00",x"01",x"01",x"02", -- 0x1EA8
		x"02",x"02",x"02",x"00",x"00",x"00",x"01",x"01", -- 0x1EB0
		x"02",x"02",x"02",x"00",x"00",x"00",x"00",x"01", -- 0x1EB8
		x"01",x"02",x"02",x"00",x"00",x"00",x"00",x"01", -- 0x1EC0
		x"01",x"02",x"02",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
		x"01",x"01",x"02",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
		x"01",x"01",x"02",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
		x"01",x"01",x"02",x"E9",x"9E",x"32",x"9F",x"7B", -- 0x1EE0
		x"9F",x"02",x"03",x"FF",x"01",x"02",x"FE",x"01", -- 0x1EE8
		x"03",x"FF",x"03",x"02",x"FE",x"01",x"02",x"FF", -- 0x1EF0
		x"02",x"02",x"FE",x"01",x"01",x"FE",x"01",x"02", -- 0x1EF8
		x"FE",x"01",x"01",x"FD",x"02",x"02",x"FE",x"01", -- 0x1F00
		x"01",x"FD",x"01",x"02",x"FE",x"01",x"01",x"FD", -- 0x1F08
		x"01",x"02",x"FE",x"01",x"01",x"FD",x"02",x"01", -- 0x1F10
		x"FE",x"02",x"01",x"FD",x"01",x"02",x"FE",x"03", -- 0x1F18
		x"01",x"FD",x"01",x"01",x"FE",x"02",x"01",x"FD", -- 0x1F20
		x"01",x"02",x"FE",x"02",x"01",x"FD",x"01",x"01", -- 0x1F28
		x"FE",x"00",x"01",x"03",x"00",x"02",x"03",x"FF", -- 0x1F30
		x"01",x"02",x"FF",x"01",x"03",x"FF",x"01",x"02", -- 0x1F38
		x"FF",x"01",x"02",x"FE",x"02",x"03",x"FF",x"01", -- 0x1F40
		x"02",x"FE",x"01",x"03",x"FF",x"02",x"02",x"FE", -- 0x1F48
		x"01",x"03",x"FF",x"09",x"02",x"FE",x"01",x"01", -- 0x1F50
		x"FE",x"02",x"02",x"FE",x"01",x"01",x"FD",x"02", -- 0x1F58
		x"02",x"FE",x"01",x"01",x"FD",x"01",x"02",x"FE", -- 0x1F60
		x"01",x"01",x"FD",x"01",x"02",x"FE",x"02",x"01", -- 0x1F68
		x"FD",x"01",x"02",x"FE",x"01",x"01",x"FD",x"01", -- 0x1F70
		x"01",x"FE",x"00",x"02",x"03",x"00",x"04",x"03", -- 0x1F78
		x"FF",x"01",x"02",x"FE",x"0B",x"03",x"FF",x"01", -- 0x1F80
		x"02",x"FE",x"01",x"03",x"FF",x"01",x"02",x"FF", -- 0x1F88
		x"01",x"02",x"FE",x"03",x"02",x"FF",x"02",x"02", -- 0x1F90
		x"FE",x"01",x"02",x"FF",x"04",x"02",x"FE",x"01", -- 0x1F98
		x"02",x"FF",x"04",x"02",x"FE",x"01",x"02",x"FE", -- 0x1FA0
		x"00",x"01",x"0C",x"00",x"01",x"05",x"0C",x"00", -- 0x1FA8
		x"00",x"01",x"0C",x"00",x"01",x"05",x"0C",x"00", -- 0x1FB0
		x"00",x"01",x"0C",x"00",x"01",x"04",x"0C",x"00", -- 0x1FB8
		x"00",x"01",x"0C",x"00",x"01",x"04",x"0C",x"00", -- 0x1FC0
		x"00",x"01",x"0C",x"00",x"01",x"04",x"0C",x"00", -- 0x1FC8
		x"00",x"01",x"0C",x"00",x"01",x"03",x"0C",x"00", -- 0x1FD0
		x"00",x"01",x"0C",x"00",x"01",x"03",x"0C",x"00", -- 0x1FD8
		x"00",x"01",x"0C",x"00",x"01",x"03",x"0C",x"00", -- 0x1FE0
		x"00",x"01",x"0C",x"00",x"01",x"03",x"0C",x"00", -- 0x1FE8
		x"00",x"01",x"0C",x"00",x"01",x"03",x"0C",x"00", -- 0x1FF0
		x"00",x"01",x"0C",x"00",x"01",x"03",x"0C",x"00", -- 0x1FF8
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2000
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2008
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2010
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2018
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2020
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2028
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2030
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2038
		x"00",x"01",x"0C",x"00",x"01",x"02",x"0C",x"00", -- 0x2040
		x"00",x"01",x"0C",x"00",x"01",x"01",x"0D",x"00", -- 0x2048
		x"00",x"01",x"0D",x"00",x"01",x"01",x"0D",x"00", -- 0x2050
		x"00",x"01",x"0D",x"00",x"01",x"01",x"0D",x"00", -- 0x2058
		x"00",x"01",x"0D",x"01",x"01",x"01",x"0D",x"00", -- 0x2060
		x"00",x"01",x"0E",x"01",x"01",x"01",x"0E",x"00", -- 0x2068
		x"00",x"01",x"0E",x"00",x"01",x"01",x"0E",x"00", -- 0x2070
		x"00",x"01",x"0E",x"01",x"01",x"01",x"0E",x"00", -- 0x2078
		x"00",x"01",x"0E",x"01",x"01",x"01",x"0E",x"00", -- 0x2080
		x"00",x"01",x"0E",x"01",x"00",x"01",x"0E",x"00", -- 0x2088
		x"00",x"01",x"0F",x"01",x"01",x"01",x"0F",x"00", -- 0x2090
		x"00",x"01",x"0F",x"01",x"01",x"01",x"0F",x"00", -- 0x2098
		x"00",x"01",x"0F",x"01",x"00",x"01",x"0F",x"00", -- 0x20A0
		x"00",x"01",x"0F",x"01",x"00",x"01",x"0F",x"00", -- 0x20A8
		x"00",x"01",x"0F",x"01",x"01",x"01",x"00",x"00", -- 0x20B0
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20B8
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20C0
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20C8
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20D0
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20D8
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20E0
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20E8
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20F0
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x20F8
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x2100
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x2108
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x2110
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x2118
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x2120
		x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00", -- 0x2128
		x"00",x"18",x"00",x"01",x"00",x"30",x"00",x"02", -- 0x2130
		x"00",x"63",x"00",x"03",x"00",x"00",x"01",x"02", -- 0x2138
		x"00",x"01",x"02",x"01",x"01",x"02",x"00",x"01", -- 0x2140
		x"02",x"01",x"01",x"02",x"00",x"07",x"02",x"01", -- 0x2148
		x"01",x"02",x"02",x"01",x"02",x"01",x"01",x"02", -- 0x2150
		x"02",x"01",x"02",x"01",x"04",x"02",x"02",x"01", -- 0x2158
		x"01",x"02",x"07",x"02",x"02",x"01",x"00",x"02", -- 0x2160
		x"01",x"01",x"02",x"01",x"00",x"02",x"01",x"01", -- 0x2168
		x"02",x"01",x"00",x"02",x"01",x"01",x"02",x"06", -- 0x2170
		x"00",x"02",x"06",x"00",x"02",x"01",x"FF",x"02", -- 0x2178
		x"01",x"00",x"02",x"01",x"FF",x"02",x"01",x"00", -- 0x2180
		x"02",x"01",x"FF",x"02",x"01",x"00",x"02",x"07", -- 0x2188
		x"FE",x"02",x"01",x"FF",x"02",x"04",x"FE",x"02", -- 0x2190
		x"01",x"FE",x"01",x"01",x"FE",x"02",x"01",x"FE", -- 0x2198
		x"01",x"01",x"FE",x"02",x"07",x"FE",x"01",x"01", -- 0x21A0
		x"FE",x"00",x"01",x"FE",x"01",x"01",x"FE",x"00", -- 0x21A8
		x"01",x"FE",x"01",x"01",x"FE",x"00",x"00",x"01", -- 0x21B0
		x"1C",x"40",x"D4",x"00",x"04",x"1C",x"41",x"D4", -- 0x21B8
		x"19",x"0B",x"1C",x"45",x"D4",x"16",x"01",x"1C", -- 0x21C0
		x"5F",x"D4",x"19",x"01",x"0A",x"7F",x"D5",x"1A", -- 0x21C8
		x"01",x"1C",x"5E",x"D4",x"33",x"06",x"17",x"90", -- 0x21D0
		x"D4",x"B0",x"01",x"1C",x"4A",x"D4",x"1A",x"00", -- 0x21D8
		x"01",x"1C",x"40",x"D4",x"00",x"1D",x"1C",x"41", -- 0x21E0
		x"D4",x"19",x"01",x"1C",x"5F",x"D4",x"19",x"01", -- 0x21E8
		x"0A",x"7F",x"D5",x"1A",x"01",x"1C",x"5E",x"D4", -- 0x21F0
		x"33",x"06",x"17",x"90",x"D4",x"B0",x"00",x"01", -- 0x21F8
		x"1C",x"4A",x"D4",x"1A",x"00",x"10",x"1C",x"41", -- 0x2200
		x"D4",x"19",x"05",x"1C",x"52",x"D4",x"10",x"01", -- 0x2208
		x"0E",x"34",x"D5",x"16",x"05",x"1C",x"4C",x"D4", -- 0x2210
		x"1A",x"00",x"1E",x"1C",x"40",x"D4",x"00",x"01", -- 0x2218
		x"1C",x"5F",x"D4",x"19",x"01",x"0A",x"7F",x"D5", -- 0x2220
		x"1A",x"01",x"1C",x"5E",x"D4",x"33",x"06",x"17", -- 0x2228
		x"90",x"D4",x"B0",x"0C",x"08",x"00",x"D5",x"1A", -- 0x2230
		x"0C",x"06",x"40",x"D4",x"19",x"0C",x"04",x"40", -- 0x2238
		x"D7",x"16",x"00",x"01",x"1C",x"59",x"D4",x"19", -- 0x2240
		x"01",x"1C",x"54",x"D4",x"16",x"01",x"1C",x"51", -- 0x2248
		x"D4",x"1A",x"01",x"1C",x"4A",x"D4",x"16",x"00", -- 0x2250
		x"1C",x"1C",x"42",x"D4",x"19",x"01",x"03",x"B4", -- 0x2258
		x"D6",x"1A",x"03",x"05",x"8A",x"D5",x"1A",x"01", -- 0x2260
		x"1C",x"4E",x"D4",x"16",x"01",x"1C",x"49",x"D4", -- 0x2268
		x"19",x"01",x"01",x"29",x"D5",x"05",x"01",x"04", -- 0x2270
		x"09",x"D6",x"1A",x"00",x"1D",x"1C",x"41",x"D4", -- 0x2278
		x"16",x"01",x"06",x"45",x"D4",x"11",x"01",x"16", -- 0x2280
		x"05",x"D5",x"13",x"01",x"12",x"48",x"D4",x"1C", -- 0x2288
		x"01",x"0A",x"88",x"D6",x"19",x"01",x"1C",x"52", -- 0x2290
		x"D4",x"1A",x"01",x"06",x"00",x"D7",x"05",x"00", -- 0x2298
		x"01",x"1C",x"5B",x"D4",x"16",x"12",x"1C",x"48", -- 0x22A0
		x"D4",x"19",x"0E",x"08",x"6C",x"D6",x"1A",x"0E", -- 0x22A8
		x"01",x"48",x"D7",x"19",x"01",x"06",x"00",x"D7", -- 0x22B0
		x"05",x"00",x"1E",x"1C",x"40",x"D4",x"00",x"01", -- 0x22B8
		x"1C",x"5F",x"D4",x"19",x"01",x"0A",x"7F",x"D5", -- 0x22C0
		x"1A",x"01",x"1C",x"5E",x"D4",x"33",x"14",x"1C", -- 0x22C8
		x"48",x"D4",x"19",x"01",x"0D",x"55",x"D5",x"1A", -- 0x22D0
		x"01",x"0E",x"32",x"D6",x"16",x"01",x"0C",x"F0", -- 0x22D8
		x"D5",x"16",x"01",x"1C",x"5C",x"D4",x"1A",x"02", -- 0x22E0
		x"1C",x"58",x"D4",x"06",x"00",x"1E",x"1C",x"40", -- 0x22E8
		x"D4",x"00",x"01",x"1C",x"5F",x"D4",x"19",x"01", -- 0x22F0
		x"0A",x"7F",x"D5",x"1A",x"01",x"1C",x"5E",x"D4", -- 0x22F8
		x"33",x"01",x"1C",x"4F",x"D4",x"16",x"0C",x"08", -- 0x2300
		x"00",x"D5",x"1A",x"0C",x"06",x"40",x"D4",x"19", -- 0x2308
		x"0C",x"04",x"40",x"D7",x"16",x"00",x"1E",x"1C", -- 0x2310
		x"40",x"D4",x"00",x"01",x"1C",x"5F",x"D4",x"19", -- 0x2318
		x"01",x"0A",x"7F",x"D5",x"1A",x"01",x"1C",x"5E", -- 0x2320
		x"D4",x"33",x"06",x"17",x"92",x"D4",x"B0",x"01", -- 0x2328
		x"1C",x"4F",x"D4",x"16",x"0C",x"08",x"00",x"D5", -- 0x2330
		x"1A",x"0C",x"06",x"40",x"D4",x"19",x"0C",x"04", -- 0x2338
		x"40",x"D7",x"16",x"00",x"30",x"30",x"30",x"30", -- 0x2340
		x"00",x"30",x"01",x"02",x"03",x"04",x"05",x"06", -- 0x2348
		x"07",x"08",x"09",x"0A",x"0B",x"0C",x"07",x"0D", -- 0x2350
		x"0E",x"0E",x"0E",x"0F",x"10",x"11",x"12",x"13", -- 0x2358
		x"13",x"14",x"15",x"16",x"17",x"16",x"18",x"30", -- 0x2360
		x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"07",x"1F", -- 0x2368
		x"20",x"21",x"22",x"23",x"07",x"24",x"25",x"26", -- 0x2370
		x"27",x"28",x"29",x"08",x"2A",x"08",x"2B",x"2C", -- 0x2378
		x"2D",x"2E",x"2F",x"2F",x"34",x"35",x"30",x"36", -- 0x2380
		x"37",x"38",x"30",x"30",x"30",x"39",x"3A",x"3B", -- 0x2388
		x"3C",x"3D",x"3E",x"3F",x"40",x"41",x"42",x"43", -- 0x2390
		x"07",x"44",x"45",x"46",x"47",x"28",x"07",x"48", -- 0x2398
		x"49",x"4A",x"4A",x"4B",x"4C",x"4D",x"4E",x"4F", -- 0x23A0
		x"50",x"51",x"52",x"53",x"54",x"55",x"56",x"57", -- 0x23A8
		x"58",x"59",x"5A",x"5B",x"5C",x"5D",x"07",x"5E", -- 0x23B0
		x"08",x"5F",x"60",x"28",x"07",x"61",x"62",x"63", -- 0x23B8
		x"64",x"28",x"07",x"08",x"65",x"66",x"67",x"2C", -- 0x23C0
		x"69",x"6A",x"6B",x"6C",x"6D",x"35",x"00",x"04", -- 0x23C8
		x"00",x"00",x"38",x"30",x"0C",x"0A",x"19",x"0C", -- 0x23D0
		x"18",x"16",x"00",x"03",x"50",x"00",x"0A",x"15", -- 0x23D8
		x"15",x"30",x"30",x"30",x"30",x"30",x"00",x"03", -- 0x23E0
		x"00",x"00",x"1B",x"12",x"10",x"11",x"1D",x"30", -- 0x23E8
		x"30",x"30",x"00",x"02",x"50",x"00",x"1B",x"0E", -- 0x23F0
		x"1C",x"0E",x"1B",x"1F",x"0E",x"0D",x"00",x"02", -- 0x23F8
		x"00",x"00",x"0E",x"21",x"0E",x"0D",x"0E",x"21", -- 0x2400
		x"0E",x"1C",x"00",x"00",x"99",x"99",x"1F",x"1E", -- 0x2408
		x"15",x"10",x"1E",x"1C",x"30",x"30",x"00",x"00", -- 0x2410
		x"88",x"88",x"1C",x"18",x"17",x"1C",x"18",x"17", -- 0x2418
		x"30",x"30",x"00",x"00",x"77",x"77",x"11",x"12", -- 0x2420
		x"10",x"0E",x"16",x"0A",x"1B",x"1E",x"00",x"00", -- 0x2428
		x"66",x"66",x"0E",x"21",x"0E",x"0D",x"0E",x"21", -- 0x2430
		x"0E",x"1C",x"00",x"00",x"55",x"55",x"17",x"0A", -- 0x2438
		x"14",x"0A",x"1C",x"0A",x"1D",x"18",x"00",x"0D", -- 0x2440
		x"22",x"D1",x"38",x"30",x"01",x"09",x"08",x"04", -- 0x2448
		x"30",x"0C",x"0A",x"19",x"0C",x"18",x"16",x"00", -- 0x2450
		x"00",x"11",x"EB",x"D0",x"19",x"1E",x"1C",x"11", -- 0x2458
		x"30",x"1C",x"1D",x"0A",x"1B",x"1D",x"30",x"0B", -- 0x2460
		x"1E",x"1D",x"1D",x"18",x"17",x"00",x"0F",x"09", -- 0x2468
		x"D1",x"18",x"17",x"0E",x"30",x"19",x"15",x"0A", -- 0x2470
		x"22",x"0E",x"1B",x"30",x"18",x"17",x"15",x"22", -- 0x2478
		x"00",x"12",x"E9",x"D0",x"18",x"17",x"0E",x"30", -- 0x2480
		x"18",x"1B",x"30",x"1D",x"20",x"18",x"30",x"19", -- 0x2488
		x"15",x"0A",x"22",x"0E",x"1B",x"1C",x"00",x"0B", -- 0x2490
		x"4A",x"D1",x"12",x"17",x"1C",x"0E",x"1B",x"1D", -- 0x2498
		x"30",x"0C",x"18",x"12",x"17",x"00",x"08",x"8B", -- 0x24A0
		x"D1",x"19",x"15",x"0A",x"22",x"0E",x"1B",x"30", -- 0x24A8
		x"01",x"00",x"08",x"8B",x"D1",x"19",x"15",x"0A", -- 0x24B0
		x"22",x"0E",x"1B",x"30",x"02",x"00",x"05",x"AD", -- 0x24B8
		x"D1",x"1B",x"0E",x"0A",x"0D",x"22",x"00",x"03", -- 0x24C0
		x"9F",x"D0",x"01",x"1E",x"19",x"0A",x"7F",x"D1", -- 0x24C8
		x"11",x"12",x"10",x"11",x"30",x"1C",x"0C",x"18", -- 0x24D0
		x"1B",x"0E",x"03",x"3F",x"D3",x"02",x"1E",x"19", -- 0x24D8
		x"00",x"06",x"A0",x"D2",x"0C",x"1B",x"0E",x"0D", -- 0x24E0
		x"12",x"1D",x"00",x"15",x"CF",x"D0",x"1D",x"18", -- 0x24E8
		x"19",x"30",x"05",x"30",x"1B",x"0A",x"17",x"14", -- 0x24F0
		x"12",x"17",x"10",x"30",x"1C",x"0C",x"18",x"1B", -- 0x24F8
		x"0E",x"28",x"28",x"03",x"8B",x"D0",x"1D",x"18", -- 0x2500
		x"19",x"03",x"88",x"D0",x"02",x"17",x"0D",x"03", -- 0x2508
		x"86",x"D0",x"03",x"1B",x"0D",x"03",x"84",x"D0", -- 0x2510
		x"04",x"1D",x"11",x"03",x"82",x"D0",x"05",x"1D", -- 0x2518
		x"11",x"00",x"16",x"AD",x"D0",x"2A",x"30",x"22", -- 0x2520
		x"18",x"1E",x"1B",x"30",x"1B",x"0A",x"17",x"14", -- 0x2528
		x"12",x"17",x"10",x"30",x"1C",x"0C",x"18",x"1B", -- 0x2530
		x"0E",x"30",x"2B",x"00",x"01",x"AD",x"D0",x"30", -- 0x2538
		x"00",x"01",x"AD",x"D0",x"30",x"00",x"09",x"6B", -- 0x2540
		x"D1",x"10",x"0A",x"16",x"0E",x"30",x"18",x"1F", -- 0x2548
		x"0E",x"1B",x"00",x"05",x"BB",x"D1",x"1D",x"12", -- 0x2550
		x"16",x"0E",x"1B",x"0F",x"35",x"D1",x"48",x"0C", -- 0x2558
		x"18",x"17",x"1D",x"12",x"17",x"1E",x"0E",x"30", -- 0x2560
		x"10",x"0A",x"16",x"0E",x"49",x"19",x"72",x"D0", -- 0x2568
		x"19",x"1E",x"1C",x"11",x"30",x"0A",x"17",x"0D", -- 0x2570
		x"30",x"11",x"18",x"15",x"0D",x"30",x"0F",x"12", -- 0x2578
		x"1B",x"0E",x"30",x"0B",x"1E",x"1D",x"1D",x"18", -- 0x2580
		x"17",x"16",x"B0",x"D0",x"1D",x"11",x"0E",x"17", -- 0x2588
		x"30",x"19",x"1E",x"1C",x"11",x"30",x"1C",x"1D", -- 0x2590
		x"0A",x"1B",x"1D",x"30",x"0B",x"1E",x"1D",x"1D", -- 0x2598
		x"18",x"17",x"19",x"6E",x"D0",x"0B",x"0E",x"0F", -- 0x25A0
		x"18",x"1B",x"0E",x"30",x"1D",x"12",x"16",x"0E", -- 0x25A8
		x"30",x"0C",x"18",x"1E",x"17",x"1D",x"30",x"0E", -- 0x25B0
		x"17",x"1D",x"0E",x"1B",x"30",x"00",x"00",x"0A", -- 0x25B8
		x"0D",x"B7",x"D0",x"1C",x"11",x"18",x"18",x"1D", -- 0x25C0
		x"12",x"17",x"10",x"30",x"0D",x"18",x"20",x"17", -- 0x25C8
		x"00",x"0A",x"0D",x"F4",x"D0",x"1C",x"11",x"18", -- 0x25D0
		x"18",x"1D",x"12",x"17",x"10",x"30",x"0D",x"18", -- 0x25D8
		x"20",x"17",x"00",x"0A",x"0B",x"B1",x"D0",x"1D", -- 0x25E0
		x"18",x"0D",x"0A",x"22",x"5B",x"1C",x"30",x"1D", -- 0x25E8
		x"18",x"19",x"00",x"0A",x"0A",x"B4",x"D0",x"19", -- 0x25F0
		x"0E",x"1B",x"0C",x"0E",x"17",x"1D",x"0A",x"10", -- 0x25F8
		x"0E",x"00",x"00",x"08",x"8E",x"D1",x"17",x"18", -- 0x2600
		x"30",x"0B",x"18",x"17",x"1E",x"1C",x"00",x"0D", -- 0x2608
		x"4E",x"D1",x"1C",x"19",x"0E",x"0C",x"12",x"0A", -- 0x2610
		x"15",x"30",x"0B",x"18",x"17",x"1E",x"1C",x"09", -- 0x2618
		x"8C",x"D1",x"05",x"00",x"00",x"00",x"00",x"30", -- 0x2620
		x"19",x"1D",x"1C",x"00",x"18",x"99",x"D0",x"2A", -- 0x2628
		x"30",x"29",x"30",x"0A",x"17",x"0D",x"30",x"19", -- 0x2630
		x"18",x"12",x"17",x"1D",x"30",x"1E",x"19",x"30", -- 0x2638
		x"1C",x"1D",x"0A",x"10",x"0E",x"30",x"2B",x"00", -- 0x2640
		x"0A",x"71",x"D1",x"15",x"0A",x"1C",x"1D",x"30", -- 0x2648
		x"1C",x"1D",x"0A",x"10",x"0E",x"00",x"04",x"31", -- 0x2650
		x"D1",x"15",x"0A",x"1C",x"1D",x"00",x"05",x"31", -- 0x2658
		x"D2",x"1C",x"1D",x"0A",x"10",x"0E",x"00",x"07", -- 0x2660
		x"29",x"D1",x"68",x"37",x"01",x"00",x"00",x"00", -- 0x2668
		x"4A",x"00",x"0A",x"0E",x"3B",x"D1",x"0C",x"18", -- 0x2670
		x"17",x"10",x"1B",x"0A",x"1D",x"1E",x"15",x"0A", -- 0x2678
		x"1D",x"12",x"18",x"17",x"00",x"0A",x"0C",x"56", -- 0x2680
		x"D1",x"20",x"0E",x"30",x"10",x"12",x"1F",x"0E", -- 0x2688
		x"30",x"1E",x"19",x"30",x"28",x"00",x"0A",x"0E", -- 0x2690
		x"30",x"D1",x"01",x"00",x"34",x"00",x"00",x"00", -- 0x2698
		x"34",x"00",x"00",x"00",x"30",x"19",x"1D",x"1C", -- 0x26A0
		x"00",x"0A",x"13",x"E8",x"D0",x"19",x"1B",x"0E", -- 0x26A8
		x"1C",x"0E",x"17",x"1D",x"0E",x"0D",x"30",x"0B", -- 0x26B0
		x"22",x"30",x"0C",x"0A",x"19",x"0C",x"18",x"16", -- 0x26B8
		x"00",x"0A",x"17",x"A5",x"D0",x"19",x"1C",x"24", -- 0x26C0
		x"30",x"11",x"18",x"19",x"0E",x"30",x"18",x"1E", -- 0x26C8
		x"1B",x"30",x"17",x"0E",x"21",x"1D",x"30",x"10", -- 0x26D0
		x"0A",x"16",x"0E",x"24",x"00",x"07",x"8F",x"D1", -- 0x26D8
		x"22",x"18",x"1E",x"30",x"0A",x"1B",x"0E",x"14", -- 0x26E0
		x"CD",x"D0",x"1D",x"11",x"0E",x"30",x"0B",x"0E", -- 0x26E8
		x"1C",x"1D",x"30",x"18",x"0F",x"30",x"19",x"15", -- 0x26F0
		x"0A",x"22",x"0E",x"1B",x"30",x"28",x"00",x"14", -- 0x26F8
		x"C8",x"D0",x"0F",x"12",x"10",x"11",x"1D",x"30", -- 0x2700
		x"15",x"0A",x"1C",x"1D",x"30",x"18",x"17",x"0E", -- 0x2708
		x"30",x"1C",x"1D",x"0A",x"10",x"0E",x"00",x"27", -- 0x2710
		x"A7",x"32",x"A7",x"3F",x"A7",x"48",x"A7",x"53", -- 0x2718
		x"A7",x"5D",x"A7",x"68",x"A7",x"74",x"A7",x"00", -- 0x2720
		x"06",x"B4",x"D1",x"16",x"12",x"0D",x"20",x"0A", -- 0x2728
		x"22",x"00",x"00",x"08",x"94",x"D1",x"16",x"0A", -- 0x2730
		x"1B",x"1C",x"11",x"0A",x"15",x"15",x"00",x"00", -- 0x2738
		x"04",x"D4",x"D1",x"0A",x"1D",x"1D",x"1E",x"00", -- 0x2740
		x"00",x"06",x"B4",x"D1",x"1B",x"0A",x"0B",x"0A", -- 0x2748
		x"1E",x"15",x"00",x"00",x"05",x"D4",x"D1",x"15", -- 0x2750
		x"0E",x"22",x"1D",x"0E",x"00",x"00",x"06",x"B4", -- 0x2758
		x"D1",x"1C",x"0A",x"12",x"19",x"0A",x"17",x"00", -- 0x2760
		x"00",x"07",x"94",x"D1",x"12",x"20",x"18",x"13", -- 0x2768
		x"12",x"16",x"0A",x"00",x"00",x"07",x"94",x"D1", -- 0x2770
		x"18",x"14",x"12",x"17",x"0A",x"20",x"0A",x"00", -- 0x2778
		x"C4",x"A7",x"C6",x"A7",x"C8",x"A7",x"CA",x"A7", -- 0x2780
		x"CC",x"A7",x"CE",x"A7",x"CF",x"A7",x"CF",x"A7", -- 0x2788
		x"CF",x"A7",x"CF",x"A7",x"CF",x"A7",x"CF",x"A7", -- 0x2790
		x"CF",x"A7",x"CF",x"A7",x"CF",x"A7",x"CF",x"A7", -- 0x2798
		x"D0",x"A7",x"D3",x"A7",x"D6",x"A7",x"D9",x"A7", -- 0x27A0
		x"DC",x"A7",x"E0",x"A7",x"E4",x"A7",x"E8",x"A7", -- 0x27A8
		x"EC",x"A7",x"EF",x"A7",x"F2",x"A7",x"F6",x"A7", -- 0x27B0
		x"FA",x"A7",x"FE",x"A7",x"02",x"A8",x"06",x"A8", -- 0x27B8
		x"0A",x"A8",x"0D",x"A8",x"00",x"FF",x"01",x"FF", -- 0x27C0
		x"02",x"FF",x"03",x"FF",x"04",x"FF",x"05",x"FF", -- 0x27C8
		x"03",x"04",x"FF",x"04",x"03",x"FF",x"03",x"03", -- 0x27D0
		x"FF",x"04",x"04",x"FF",x"03",x"03",x"04",x"FF", -- 0x27D8
		x"04",x"04",x"03",x"FF",x"03",x"04",x"03",x"FF", -- 0x27E0
		x"04",x"03",x"04",x"FF",x"03",x"01",x"FF",x"04", -- 0x27E8
		x"01",x"FF",x"00",x"00",x"01",x"FF",x"00",x"00", -- 0x27F0
		x"02",x"FF",x"00",x"00",x"03",x"FF",x"00",x"00", -- 0x27F8
		x"04",x"FF",x"00",x"05",x"03",x"FF",x"00",x"05", -- 0x2800
		x"04",x"FF",x"05",x"03",x"FF",x"05",x"04",x"FF", -- 0x2808
		x"3F",x"60",x"3F",x"C0",x"7C",x"A8",x"5C",x"A8", -- 0x2810
		x"3C",x"A8",x"1C",x"A8",x"40",x"40",x"30",x"40", -- 0x2818
		x"30",x"30",x"30",x"40",x"30",x"30",x"30",x"40", -- 0x2820
		x"30",x"20",x"20",x"40",x"30",x"20",x"20",x"40", -- 0x2828
		x"20",x"20",x"20",x"40",x"20",x"20",x"20",x"40", -- 0x2830
		x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40", -- 0x2838
		x"40",x"30",x"30",x"40",x"40",x"40",x"30",x"40", -- 0x2840
		x"30",x"30",x"20",x"40",x"40",x"40",x"30",x"40", -- 0x2848
		x"30",x"30",x"30",x"40",x"30",x"30",x"30",x"40", -- 0x2850
		x"30",x"30",x"30",x"40",x"30",x"30",x"20",x"30", -- 0x2858
		x"20",x"20",x"20",x"30",x"20",x"20",x"10",x"20", -- 0x2860
		x"20",x"10",x"10",x"20",x"20",x"10",x"10",x"20", -- 0x2868
		x"10",x"10",x"10",x"20",x"10",x"10",x"10",x"20", -- 0x2870
		x"10",x"10",x"10",x"30",x"30",x"20",x"20",x"20", -- 0x2878
		x"20",x"10",x"10",x"10",x"10",x"10",x"10",x"10", -- 0x2880
		x"10",x"10",x"10",x"10",x"30",x"20",x"10",x"10", -- 0x2888
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10", -- 0x2890
		x"10",x"10",x"10",x"20",x"B0",x"A8",x"AC",x"A8", -- 0x2898
		x"A4",x"A8",x"A8",x"A8",x"80",x"70",x"60",x"50", -- 0x28A0
		x"80",x"60",x"40",x"30",x"40",x"40",x"30",x"30", -- 0x28A8
		x"40",x"30",x"30",x"30",x"07",x"04",x"40",x"00", -- 0x28B0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28B8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28C0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28C8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28D0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28D8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28E0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28E8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28F0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x28F8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2900
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2908
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2910
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2918
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2920
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2928
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2930
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2938
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2940
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2948
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2950
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2958
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2960
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2968
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2970
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2978
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2980
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2988
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2990
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2998
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29A0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29A8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29B0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29B8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29C0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29C8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29D0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29D8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29E0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29E8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29F0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x29F8
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A00
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A08
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A10
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A18
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A20
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A28
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A30
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A38
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A40
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A48
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A50
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A58
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A60
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A68
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A70
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A78
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A80
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A88
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A90
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2A98
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2AA0
		x"07",x"04",x"40",x"00",x"07",x"04",x"40",x"00", -- 0x2AA8
		x"07",x"04",x"40",x"00",x"C4",x"AA",x"29",x"AB", -- 0x2AB0
		x"97",x"AB",x"46",x"AC",x"61",x"AD",x"E3",x"AD", -- 0x2AB8
		x"90",x"AE",x"D5",x"AF",x"4D",x"0C",x"00",x"02", -- 0x2AC0
		x"01",x"0D",x"01",x"02",x"01",x"0D",x"00",x"02", -- 0x2AC8
		x"04",x"0D",x"01",x"02",x"09",x"0E",x"01",x"01", -- 0x2AD0
		x"01",x"0E",x"02",x"00",x"01",x"0F",x"01",x"01", -- 0x2AD8
		x"01",x"0F",x"02",x"00",x"34",x"00",x"02",x"00", -- 0x2AE0
		x"01",x"01",x"02",x"00",x"01",x"01",x"01",x"FF", -- 0x2AE8
		x"01",x"02",x"02",x"00",x"09",x"02",x"01",x"FF", -- 0x2AF0
		x"04",x"03",x"01",x"FE",x"01",x"03",x"00",x"FE", -- 0x2AF8
		x"01",x"03",x"01",x"FE",x"0E",x"04",x"00",x"FE", -- 0x2B00
		x"01",x"05",x"FF",x"FE",x"01",x"05",x"00",x"FE", -- 0x2B08
		x"04",x"05",x"FF",x"FE",x"09",x"06",x"FF",x"FF", -- 0x2B10
		x"01",x"06",x"FE",x"00",x"01",x"07",x"FF",x"FF", -- 0x2B18
		x"01",x"07",x"FE",x"00",x"63",x"08",x"FE",x"00", -- 0x2B20
		x"00",x"64",x"08",x"FE",x"00",x"02",x"09",x"FE", -- 0x2B28
		x"00",x"05",x"09",x"FE",x"01",x"01",x"0A",x"FE", -- 0x2B30
		x"02",x"01",x"0A",x"FF",x"02",x"01",x"0A",x"FE", -- 0x2B38
		x"02",x"04",x"0B",x"FF",x"02",x"01",x"0B",x"00", -- 0x2B40
		x"02",x"01",x"0B",x"FF",x"02",x"19",x"0C",x"00", -- 0x2B48
		x"02",x"01",x"0D",x"01",x"02",x"01",x"0D",x"00", -- 0x2B50
		x"02",x"04",x"0D",x"01",x"02",x"01",x"0E",x"02", -- 0x2B58
		x"02",x"01",x"0E",x"01",x"02",x"01",x"0E",x"02", -- 0x2B60
		x"02",x"05",x"0F",x"02",x"01",x"02",x"0F",x"02", -- 0x2B68
		x"00",x"58",x"00",x"02",x"00",x"01",x"01",x"02", -- 0x2B70
		x"FE",x"01",x"02",x"01",x"FF",x"01",x"03",x"01", -- 0x2B78
		x"FE",x"FF",x"00",x"04",x"00",x"FE",x"01",x"05", -- 0x2B80
		x"FF",x"FE",x"01",x"06",x"FF",x"FF",x"01",x"07", -- 0x2B88
		x"FE",x"FE",x"63",x"08",x"FE",x"00",x"00",x"1F", -- 0x2B90
		x"08",x"FE",x"00",x"FF",x"01",x"08",x"FE",x"00", -- 0x2B98
		x"01",x"09",x"FE",x"00",x"04",x"09",x"FE",x"01", -- 0x2BA0
		x"02",x"0A",x"FE",x"02",x"03",x"0B",x"FF",x"02", -- 0x2BA8
		x"01",x"0B",x"00",x"02",x"40",x"0C",x"00",x"02", -- 0x2BB0
		x"01",x"0D",x"00",x"02",x"03",x"0D",x"01",x"02", -- 0x2BB8
		x"02",x"0E",x"02",x"02",x"04",x"0F",x"02",x"01", -- 0x2BC0
		x"01",x"0F",x"02",x"00",x"0B",x"00",x"02",x"00", -- 0x2BC8
		x"FF",x"02",x"00",x"02",x"00",x"01",x"01",x"02", -- 0x2BD0
		x"00",x"03",x"01",x"02",x"FF",x"04",x"02",x"02", -- 0x2BD8
		x"FE",x"01",x"02",x"01",x"FE",x"01",x"02",x"01", -- 0x2BE0
		x"FF",x"04",x"02",x"01",x"FE",x"01",x"03",x"01", -- 0x2BE8
		x"FE",x"01",x"03",x"00",x"FE",x"01",x"03",x"01", -- 0x2BF0
		x"FE",x"0C",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x2BF8
		x"FE",x"01",x"04",x"00",x"FE",x"01",x"04",x"FF", -- 0x2C00
		x"FE",x"04",x"05",x"FF",x"FE",x"01",x"05",x"FF", -- 0x2C08
		x"FF",x"01",x"05",x"FF",x"FE",x"04",x"06",x"FE", -- 0x2C10
		x"FE",x"03",x"07",x"FE",x"FF",x"01",x"07",x"FE", -- 0x2C18
		x"00",x"44",x"40",x"FE",x"00",x"06",x"41",x"FE", -- 0x2C20
		x"00",x"04",x"42",x"FE",x"00",x"04",x"42",x"FF", -- 0x2C28
		x"00",x"05",x"42",x"00",x"00",x"04",x"42",x"01", -- 0x2C30
		x"00",x"04",x"42",x"02",x"00",x"06",x"43",x"02", -- 0x2C38
		x"00",x"C7",x"44",x"02",x"00",x"00",x"1B",x"08", -- 0x2C40
		x"FE",x"00",x"FF",x"03",x"08",x"FE",x"00",x"02", -- 0x2C48
		x"09",x"FE",x"01",x"02",x"0A",x"FE",x"01",x"01", -- 0x2C50
		x"0A",x"FE",x"02",x"03",x"0A",x"FF",x"02",x"01", -- 0x2C58
		x"0B",x"FF",x"02",x"01",x"0B",x"00",x"02",x"46", -- 0x2C60
		x"0C",x"00",x"02",x"01",x"0D",x"00",x"02",x"01", -- 0x2C68
		x"0D",x"01",x"02",x"03",x"0E",x"01",x"02",x"01", -- 0x2C70
		x"0E",x"02",x"02",x"02",x"0E",x"02",x"01",x"02", -- 0x2C78
		x"0F",x"02",x"01",x"0F",x"00",x"02",x"00",x"FF", -- 0x2C80
		x"04",x"00",x"02",x"00",x"01",x"01",x"02",x"00", -- 0x2C88
		x"03",x"01",x"02",x"FF",x"02",x"02",x"02",x"FE", -- 0x2C90
		x"02",x"02",x"01",x"FE",x"01",x"02",x"01",x"FE", -- 0x2C98
		x"01",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x2CA0
		x"01",x"03",x"00",x"FE",x"02",x"04",x"00",x"FE", -- 0x2CA8
		x"01",x"05",x"00",x"FE",x"01",x"05",x"FF",x"FE", -- 0x2CB0
		x"01",x"05",x"00",x"FE",x"01",x"06",x"FF",x"FE", -- 0x2CB8
		x"02",x"06",x"FF",x"FE",x"02",x"06",x"FE",x"FE", -- 0x2CC0
		x"03",x"07",x"FE",x"FF",x"01",x"07",x"FE",x"00", -- 0x2CC8
		x"10",x"20",x"FE",x"00",x"01",x"21",x"FE",x"FF", -- 0x2CD0
		x"01",x"21",x"FE",x"00",x"02",x"21",x"FE",x"FF", -- 0x2CD8
		x"01",x"21",x"FE",x"00",x"0A",x"21",x"FE",x"FF", -- 0x2CE0
		x"01",x"21",x"FE",x"00",x"08",x"21",x"FE",x"FF", -- 0x2CE8
		x"05",x"22",x"FE",x"FF",x"01",x"22",x"FE",x"FE", -- 0x2CF0
		x"02",x"22",x"FE",x"FF",x"01",x"22",x"FE",x"FE", -- 0x2CF8
		x"01",x"22",x"FE",x"FF",x"03",x"22",x"FE",x"FE", -- 0x2D00
		x"02",x"22",x"FE",x"FF",x"02",x"22",x"FE",x"FE", -- 0x2D08
		x"02",x"22",x"FE",x"FF",x"02",x"22",x"FE",x"FE", -- 0x2D10
		x"02",x"22",x"FE",x"FF",x"02",x"22",x"FE",x"FE", -- 0x2D18
		x"02",x"22",x"FE",x"FF",x"02",x"23",x"FE",x"FE", -- 0x2D20
		x"02",x"23",x"FE",x"FF",x"03",x"23",x"FE",x"FE", -- 0x2D28
		x"01",x"23",x"FE",x"FF",x"01",x"23",x"FE",x"FE", -- 0x2D30
		x"01",x"23",x"FE",x"FF",x"01",x"23",x"FE",x"FE", -- 0x2D38
		x"01",x"23",x"FE",x"FF",x"03",x"23",x"FE",x"FE", -- 0x2D40
		x"01",x"23",x"FE",x"FF",x"05",x"23",x"FE",x"FE", -- 0x2D48
		x"01",x"23",x"FE",x"FF",x"06",x"23",x"FE",x"FE", -- 0x2D50
		x"01",x"23",x"FF",x"FE",x"63",x"23",x"FE",x"FE", -- 0x2D58
		x"00",x"28",x"0C",x"00",x"02",x"03",x"0D",x"00", -- 0x2D60
		x"02",x"03",x"0D",x"01",x"03",x"01",x"0D",x"01", -- 0x2D68
		x"02",x"01",x"0E",x"02",x"02",x"01",x"0E",x"02", -- 0x2D70
		x"01",x"01",x"0E",x"02",x"02",x"02",x"0F",x"02", -- 0x2D78
		x"01",x"01",x"0F",x"02",x"00",x"09",x"30",x"02", -- 0x2D80
		x"00",x"FF",x"05",x"30",x"02",x"00",x"06",x"31", -- 0x2D88
		x"02",x"00",x"04",x"32",x"02",x"00",x"04",x"32", -- 0x2D90
		x"01",x"00",x"05",x"32",x"00",x"00",x"04",x"32", -- 0x2D98
		x"FF",x"00",x"04",x"32",x"FE",x"00",x"06",x"33", -- 0x2DA0
		x"FE",x"00",x"06",x"34",x"FE",x"00",x"06",x"24", -- 0x2DA8
		x"FE",x"00",x"06",x"25",x"FE",x"00",x"0A",x"26", -- 0x2DB0
		x"FE",x"00",x"0C",x"27",x"FE",x"00",x"10",x"20", -- 0x2DB8
		x"FE",x"00",x"0C",x"21",x"FE",x"00",x"0A",x"22", -- 0x2DC0
		x"FE",x"00",x"06",x"23",x"FE",x"00",x"06",x"24", -- 0x2DC8
		x"FE",x"00",x"06",x"25",x"FE",x"00",x"0A",x"26", -- 0x2DD0
		x"FE",x"00",x"0C",x"27",x"FE",x"00",x"63",x"20", -- 0x2DD8
		x"FE",x"00",x"00",x"63",x"00",x"02",x"00",x"05", -- 0x2DE0
		x"0F",x"02",x"01",x"02",x"0E",x"02",x"02",x"03", -- 0x2DE8
		x"0E",x"01",x"02",x"01",x"0D",x"00",x"02",x"01", -- 0x2DF0
		x"0D",x"01",x"02",x"4E",x"0C",x"00",x"02",x"01", -- 0x2DF8
		x"0B",x"FF",x"02",x"01",x"0B",x"00",x"02",x"03", -- 0x2E00
		x"0A",x"FF",x"02",x"02",x"0A",x"FE",x"02",x"05", -- 0x2E08
		x"09",x"FE",x"01",x"06",x"08",x"FE",x"00",x"05", -- 0x2E10
		x"07",x"FE",x"FF",x"02",x"06",x"FE",x"FE",x"03", -- 0x2E18
		x"06",x"FF",x"FE",x"01",x"05",x"00",x"FE",x"01", -- 0x2E20
		x"05",x"FF",x"FE",x"4E",x"04",x"00",x"FE",x"01", -- 0x2E28
		x"05",x"FF",x"FE",x"01",x"05",x"00",x"FE",x"03", -- 0x2E30
		x"06",x"FF",x"FE",x"02",x"06",x"FE",x"FE",x"05", -- 0x2E38
		x"07",x"FE",x"FF",x"06",x"08",x"FE",x"00",x"05", -- 0x2E40
		x"09",x"FE",x"01",x"02",x"0A",x"FE",x"02",x"03", -- 0x2E48
		x"0A",x"FF",x"02",x"01",x"0B",x"00",x"02",x"01", -- 0x2E50
		x"0B",x"FF",x"02",x"4E",x"0C",x"00",x"02",x"01", -- 0x2E58
		x"0B",x"FF",x"02",x"01",x"0B",x"00",x"02",x"03", -- 0x2E60
		x"0A",x"FF",x"02",x"02",x"0A",x"FE",x"02",x"05", -- 0x2E68
		x"09",x"FE",x"01",x"06",x"08",x"FE",x"00",x"05", -- 0x2E70
		x"07",x"FE",x"FF",x"02",x"06",x"FE",x"FE",x"03", -- 0x2E78
		x"06",x"FF",x"FE",x"01",x"05",x"00",x"FE",x"01", -- 0x2E80
		x"05",x"FF",x"FE",x"66",x"04",x"00",x"FE",x"00", -- 0x2E88
		x"1B",x"08",x"FE",x"00",x"01",x"09",x"FE",x"01", -- 0x2E90
		x"01",x"09",x"FE",x"00",x"03",x"09",x"FE",x"01", -- 0x2E98
		x"04",x"0A",x"FE",x"02",x"06",x"0A",x"FF",x"02", -- 0x2EA0
		x"01",x"0B",x"00",x"02",x"01",x"0B",x"FF",x"02", -- 0x2EA8
		x"02",x"0B",x"00",x"02",x"01",x"0B",x"FF",x"02", -- 0x2EB0
		x"06",x"0C",x"00",x"02",x"01",x"0D",x"01",x"02", -- 0x2EB8
		x"02",x"0D",x"00",x"02",x"01",x"0D",x"01",x"02", -- 0x2EC0
		x"01",x"0D",x"00",x"02",x"06",x"0E",x"01",x"02", -- 0x2EC8
		x"04",x"0E",x"02",x"02",x"03",x"0F",x"02",x"01", -- 0x2ED0
		x"01",x"0F",x"02",x"00",x"01",x"0F",x"02",x"01", -- 0x2ED8
		x"06",x"00",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x2EE0
		x"01",x"01",x"02",x"00",x"03",x"01",x"02",x"FF", -- 0x2EE8
		x"04",x"02",x"02",x"FE",x"06",x"02",x"01",x"FE", -- 0x2EF0
		x"01",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x2EF8
		x"02",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x2F00
		x"06",x"04",x"00",x"FE",x"01",x"05",x"FF",x"FE", -- 0x2F08
		x"02",x"05",x"00",x"FE",x"01",x"05",x"FF",x"FE", -- 0x2F10
		x"01",x"05",x"00",x"FE",x"06",x"06",x"FF",x"FE", -- 0x2F18
		x"04",x"06",x"FE",x"FE",x"03",x"07",x"FE",x"FF", -- 0x2F20
		x"01",x"07",x"FE",x"00",x"01",x"07",x"FE",x"FF", -- 0x2F28
		x"36",x"08",x"FE",x"00",x"01",x"09",x"FE",x"01", -- 0x2F30
		x"01",x"09",x"FE",x"00",x"03",x"09",x"FE",x"01", -- 0x2F38
		x"04",x"0A",x"FE",x"02",x"06",x"0A",x"FF",x"02", -- 0x2F40
		x"01",x"0B",x"00",x"02",x"01",x"0B",x"FF",x"02", -- 0x2F48
		x"02",x"0B",x"00",x"02",x"01",x"0B",x"FF",x"02", -- 0x2F50
		x"06",x"0C",x"00",x"02",x"01",x"0D",x"01",x"02", -- 0x2F58
		x"02",x"0D",x"00",x"02",x"01",x"0D",x"01",x"02", -- 0x2F60
		x"01",x"0D",x"00",x"02",x"06",x"0E",x"01",x"02", -- 0x2F68
		x"04",x"0E",x"02",x"02",x"03",x"0F",x"02",x"01", -- 0x2F70
		x"01",x"0F",x"02",x"00",x"01",x"0F",x"02",x"01", -- 0x2F78
		x"06",x"00",x"02",x"00",x"01",x"01",x"02",x"FF", -- 0x2F80
		x"01",x"01",x"02",x"00",x"03",x"01",x"02",x"FF", -- 0x2F88
		x"04",x"02",x"02",x"FE",x"06",x"02",x"01",x"FE", -- 0x2F90
		x"01",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x2F98
		x"02",x"03",x"00",x"FE",x"01",x"03",x"01",x"FE", -- 0x2FA0
		x"06",x"04",x"00",x"FE",x"01",x"05",x"FF",x"FE", -- 0x2FA8
		x"02",x"05",x"00",x"FE",x"01",x"05",x"FF",x"FE", -- 0x2FB0
		x"01",x"05",x"00",x"FE",x"06",x"06",x"FF",x"FE", -- 0x2FB8
		x"04",x"06",x"FE",x"FE",x"03",x"07",x"FE",x"FF", -- 0x2FC0
		x"01",x"07",x"FE",x"00",x"01",x"07",x"FE",x"FF", -- 0x2FC8
		x"66",x"08",x"FE",x"00",x"00",x"2B",x"0C",x"00", -- 0x2FD0
		x"02",x"01",x"28",x"FF",x"02",x"01",x"29",x"FF", -- 0x2FD8
		x"02",x"01",x"29",x"00",x"02",x"05",x"29",x"FF", -- 0x2FE0
		x"02",x"01",x"29",x"FE",x"02",x"02",x"29",x"FF", -- 0x2FE8
		x"02",x"01",x"2A",x"FE",x"02",x"01",x"2A",x"FF", -- 0x2FF0
		x"02",x"03",x"2A",x"FE",x"02",x"01",x"2A",x"FF", -- 0x2FF8
		x"02",x"01",x"2A",x"FE",x"02",x"01",x"2A",x"FF", -- 0x3000
		x"02",x"01",x"2A",x"FE",x"02",x"05",x"29",x"FF", -- 0x3008
		x"02",x"01",x"28",x"00",x"02",x"01",x"28",x"FF", -- 0x3010
		x"02",x"0C",x"48",x"00",x"02",x"06",x"49",x"00", -- 0x3018
		x"02",x"04",x"49",x"00",x"02",x"04",x"4A",x"00", -- 0x3020
		x"01",x"05",x"4B",x"00",x"00",x"04",x"4C",x"00", -- 0x3028
		x"FF",x"04",x"4C",x"00",x"FE",x"06",x"4C",x"00", -- 0x3030
		x"FE",x"C7",x"4C",x"00",x"FE",x"00",x"4E",x"B0", -- 0x3038
		x"76",x"B0",x"9E",x"B0",x"C6",x"B0",x"EE",x"B0", -- 0x3040
		x"16",x"B1",x"3E",x"B1",x"66",x"B1",x"00",x"00", -- 0x3048
		x"00",x"04",x"00",x"F0",x"88",x"04",x"00",x"00", -- 0x3050
		x"10",x"04",x"00",x"F0",x"98",x"04",x"00",x"00", -- 0x3058
		x"20",x"04",x"00",x"F0",x"A8",x"04",x"00",x"00", -- 0x3060
		x"30",x"04",x"00",x"F0",x"B8",x"04",x"00",x"00", -- 0x3068
		x"40",x"04",x"00",x"F0",x"C8",x"04",x"00",x"00", -- 0x3070
		x"00",x"14",x"00",x"C0",x"88",x"14",x"00",x"00", -- 0x3078
		x"10",x"14",x"00",x"C0",x"98",x"14",x"00",x"00", -- 0x3080
		x"20",x"14",x"00",x"C0",x"A8",x"14",x"00",x"00", -- 0x3088
		x"30",x"14",x"00",x"C0",x"B8",x"14",x"00",x"00", -- 0x3090
		x"40",x"14",x"00",x"C0",x"C8",x"14",x"00",x"00", -- 0x3098
		x"00",x"14",x"00",x"A0",x"88",x"14",x"00",x"00", -- 0x30A0
		x"10",x"14",x"00",x"A0",x"98",x"14",x"00",x"00", -- 0x30A8
		x"20",x"14",x"00",x"A0",x"A8",x"14",x"00",x"00", -- 0x30B0
		x"30",x"14",x"00",x"A0",x"B8",x"14",x"00",x"00", -- 0x30B8
		x"40",x"14",x"00",x"A0",x"C8",x"14",x"00",x"00", -- 0x30C0
		x"08",x"14",x"00",x"C0",x"80",x"14",x"00",x"00", -- 0x30C8
		x"18",x"14",x"00",x"C0",x"90",x"14",x"00",x"00", -- 0x30D0
		x"28",x"14",x"00",x"C0",x"A0",x"14",x"00",x"00", -- 0x30D8
		x"38",x"14",x"00",x"C0",x"B0",x"14",x"00",x"00", -- 0x30E0
		x"48",x"14",x"00",x"C0",x"C0",x"14",x"00",x"00", -- 0x30E8
		x"00",x"04",x"00",x"F0",x"88",x"04",x"E0",x"00", -- 0x30F0
		x"00",x"04",x"E0",x"F0",x"88",x"04",x"C0",x"00", -- 0x30F8
		x"00",x"04",x"C0",x"F0",x"88",x"04",x"A0",x"00", -- 0x3100
		x"00",x"04",x"A0",x"F0",x"88",x"04",x"80",x"00", -- 0x3108
		x"00",x"04",x"80",x"F0",x"88",x"04",x"F0",x"00", -- 0x3110
		x"00",x"14",x"F0",x"C0",x"80",x"14",x"F0",x"00", -- 0x3118
		x"10",x"14",x"F0",x"C0",x"90",x"14",x"F0",x"00", -- 0x3120
		x"20",x"14",x"F0",x"C0",x"A0",x"14",x"F0",x"00", -- 0x3128
		x"30",x"14",x"F0",x"C0",x"B0",x"14",x"F0",x"00", -- 0x3130
		x"40",x"14",x"F0",x"C0",x"C0",x"14",x"00",x"00", -- 0x3138
		x"00",x"14",x"00",x"A0",x"80",x"14",x"00",x"00", -- 0x3140
		x"10",x"14",x"00",x"A0",x"90",x"14",x"00",x"00", -- 0x3148
		x"20",x"14",x"00",x"A0",x"A0",x"14",x"00",x"00", -- 0x3150
		x"30",x"14",x"00",x"A0",x"B0",x"14",x"00",x"00", -- 0x3158
		x"40",x"14",x"00",x"A0",x"C0",x"14",x"00",x"00", -- 0x3160
		x"00",x"04",x"00",x"F0",x"80",x"04",x"E0",x"00", -- 0x3168
		x"10",x"04",x"E0",x"F0",x"90",x"04",x"C0",x"00", -- 0x3170
		x"20",x"04",x"C0",x"F0",x"A0",x"04",x"A0",x"00", -- 0x3178
		x"30",x"04",x"A0",x"F0",x"B0",x"04",x"80",x"00", -- 0x3180
		x"40",x"04",x"80",x"F0",x"C0",x"04",x"9A",x"B1", -- 0x3188
		x"A4",x"B1",x"A4",x"B1",x"AE",x"B1",x"AE",x"B1", -- 0x3190
		x"B8",x"B1",x"21",x"21",x"19",x"19",x"11",x"11", -- 0x3198
		x"09",x"09",x"01",x"01",x"49",x"41",x"39",x"31", -- 0x31A0
		x"29",x"21",x"19",x"11",x"09",x"01",x"41",x"49", -- 0x31A8
		x"31",x"39",x"21",x"29",x"11",x"19",x"01",x"09", -- 0x31B0
		x"01",x"01",x"11",x"11",x"21",x"21",x"31",x"31", -- 0x31B8
		x"41",x"41",x"0C",x"08",x"61",x"18",x"06",x"09", -- 0x31C0
		x"31",x"30",x"06",x"09",x"31",x"30",x"06",x"0A", -- 0x31C8
		x"29",x"40",x"06",x"0A",x"21",x"50",x"06",x"0B", -- 0x31D0
		x"21",x"50",x"06",x"0B",x"21",x"50",x"06",x"0B", -- 0x31D8
		x"21",x"60",x"06",x"0C",x"21",x"60",x"06",x"0C", -- 0x31E0
		x"21",x"60",x"06",x"0C",x"21",x"60",x"06",x"0C", -- 0x31E8
		x"19",x"60",x"06",x"0C",x"11",x"60",x"06",x"0C", -- 0x31F0
		x"11",x"60",x"06",x"0D",x"09",x"60",x"06",x"0D", -- 0x31F8
		x"09",x"50",x"06",x"0D",x"00",x"50",x"06",x"0E", -- 0x3200
		x"08",x"40",x"06",x"0E",x"10",x"30",x"06",x"0F", -- 0x3208
		x"18",x"30",x"06",x"00",x"20",x"20",x"06",x"00", -- 0x3210
		x"20",x"21",x"06",x"01",x"18",x"31",x"06",x"02", -- 0x3218
		x"10",x"31",x"06",x"02",x"08",x"41",x"06",x"03", -- 0x3220
		x"00",x"51",x"06",x"03",x"00",x"51",x"06",x"03", -- 0x3228
		x"00",x"61",x"06",x"04",x"00",x"61",x"06",x"04", -- 0x3230
		x"00",x"61",x"06",x"04",x"11",x"61",x"06",x"04", -- 0x3238
		x"21",x"61",x"06",x"04",x"31",x"61",x"06",x"04", -- 0x3240
		x"31",x"61",x"06",x"05",x"39",x"61",x"06",x"05", -- 0x3248
		x"39",x"51",x"06",x"05",x"41",x"51",x"06",x"06", -- 0x3250
		x"41",x"41",x"06",x"06",x"49",x"31",x"06",x"07", -- 0x3258
		x"51",x"29",x"06",x"07",x"51",x"29",x"0C",x"08", -- 0x3260
		x"61",x"19",x"00",x"7B",x"B2",x"8F",x"B2",x"A3", -- 0x3268
		x"B2",x"B7",x"B2",x"CB",x"B2",x"DF",x"B2",x"F3", -- 0x3270
		x"B2",x"07",x"B3",x"00",x"00",x"00",x"70",x"00", -- 0x3278
		x"50",x"10",x"70",x"00",x"A0",x"20",x"70",x"00", -- 0x3280
		x"28",x"08",x"70",x"00",x"78",x"18",x"70",x"00", -- 0x3288
		x"00",x"00",x"70",x"00",x"50",x"18",x"70",x"00", -- 0x3290
		x"B0",x"18",x"70",x"00",x"28",x"0C",x"70",x"00", -- 0x3298
		x"D8",x"0C",x"70",x"00",x"00",x"00",x"70",x"00", -- 0x32A0
		x"A0",x"10",x"70",x"00",x"28",x"20",x"70",x"00", -- 0x32A8
		x"50",x"08",x"70",x"00",x"78",x"18",x"70",x"00", -- 0x32B0
		x"00",x"18",x"70",x"00",x"D8",x"24",x"70",x"00", -- 0x32B8
		x"28",x"30",x"70",x"00",x"B0",x"00",x"70",x"00", -- 0x32C0
		x"50",x"0C",x"70",x"00",x"00",x"00",x"70",x"00", -- 0x32C8
		x"00",x"10",x"70",x"00",x"00",x"20",x"70",x"00", -- 0x32D0
		x"00",x"30",x"70",x"00",x"00",x"3F",x"70",x"00", -- 0x32D8
		x"00",x"00",x"70",x"00",x"80",x"10",x"70",x"00", -- 0x32E0
		x"20",x"20",x"70",x"00",x"A0",x"30",x"70",x"00", -- 0x32E8
		x"50",x"3F",x"70",x"00",x"00",x"00",x"70",x"00", -- 0x32F0
		x"78",x"10",x"70",x"00",x"3C",x"20",x"70",x"00", -- 0x32F8
		x"00",x"30",x"70",x"00",x"78",x"3F",x"70",x"00", -- 0x3300
		x"00",x"00",x"70",x"00",x"B0",x"18",x"70",x"00", -- 0x3308
		x"60",x"30",x"70",x"00",x"D8",x"0C",x"70",x"00", -- 0x3310
		x"88",x"24",x"70",x"00",x"00",x"00",x"70",x"00", -- 0x3318
		x"90",x"80",x"70",x"00",x"00",x"10",x"70",x"00", -- 0x3320
		x"90",x"90",x"70",x"00",x"00",x"20",x"70",x"00", -- 0x3328
		x"00",x"80",x"70",x"00",x"70",x"00",x"70",x"00", -- 0x3330
		x"00",x"90",x"70",x"00",x"70",x"10",x"70",x"00", -- 0x3338
		x"00",x"A0",x"70",x"B3",x"C0",x"B3",x"D4",x"B3", -- 0x3340
		x"00",x"00",x"00",x"70",x"00",x"50",x"10",x"70", -- 0x3348
		x"00",x"A0",x"20",x"70",x"00",x"28",x"08",x"70", -- 0x3350
		x"00",x"78",x"18",x"70",x"00",x"00",x"00",x"70", -- 0x3358
		x"00",x"50",x"18",x"70",x"00",x"B0",x"18",x"70", -- 0x3360
		x"00",x"28",x"0C",x"70",x"00",x"D8",x"0C",x"70", -- 0x3368
		x"00",x"00",x"00",x"70",x"00",x"A0",x"10",x"70", -- 0x3370
		x"00",x"28",x"20",x"70",x"00",x"50",x"08",x"70", -- 0x3378
		x"00",x"78",x"18",x"70",x"00",x"00",x"18",x"70", -- 0x3380
		x"00",x"D8",x"24",x"70",x"00",x"28",x"30",x"70", -- 0x3388
		x"00",x"B0",x"00",x"70",x"00",x"50",x"0C",x"70", -- 0x3390
		x"00",x"00",x"00",x"70",x"00",x"00",x"10",x"70", -- 0x3398
		x"00",x"00",x"20",x"70",x"00",x"00",x"30",x"70", -- 0x33A0
		x"00",x"00",x"3F",x"70",x"00",x"00",x"00",x"70", -- 0x33A8
		x"00",x"80",x"10",x"70",x"00",x"20",x"20",x"70", -- 0x33B0
		x"00",x"A0",x"30",x"70",x"00",x"50",x"3F",x"70", -- 0x33B8
		x"00",x"00",x"00",x"70",x"00",x"78",x"10",x"70", -- 0x33C0
		x"00",x"3C",x"20",x"70",x"00",x"00",x"30",x"70", -- 0x33C8
		x"00",x"78",x"3F",x"70",x"00",x"00",x"00",x"70", -- 0x33D0
		x"00",x"B0",x"18",x"70",x"00",x"60",x"30",x"70", -- 0x33D8
		x"00",x"D8",x"0C",x"70",x"00",x"88",x"24",x"70", -- 0x33E0
		x"00",x"00",x"00",x"70",x"00",x"90",x"80",x"70", -- 0x33E8
		x"00",x"00",x"10",x"70",x"00",x"90",x"90",x"70", -- 0x33F0
		x"00",x"00",x"20",x"70",x"00",x"00",x"80",x"70", -- 0x33F8
		x"00",x"70",x"00",x"70",x"00",x"00",x"90",x"70", -- 0x3400
		x"00",x"70",x"10",x"70",x"00",x"00",x"A0",x"70", -- 0x3408
		x"70",x"00",x"70",x"00",x"00",x"90",x"70",x"00", -- 0x3410
		x"70",x"10",x"70",x"00",x"00",x"A0",x"70",x"06", -- 0x3418
		x"48",x"1F",x"C6",x"E1",x"31",x"90",x"D0",x"20", -- 0x3420
		x"EF",x"D7",x"B3",x"88",x"98",x"29",x"F0",x"21", -- 0x3428
		x"DD",x"B4",x"A3",x"8B",x"A3",x"63",x"74",x"0C", -- 0x3430
		x"FE",x"E4",x"F5",x"B5",x"96",x"06",x"1D",x"3B", -- 0x3438
		x"9B",x"FF",x"C7",x"73",x"AA",x"9F",x"7D",x"1D", -- 0x3440
		x"EA",x"DC",x"E7",x"85",x"4A",x"08",x"34",x"CA", -- 0x3448
		x"5B",x"A9",x"81",x"C5",x"73",x"2C",x"59",x"25", -- 0x3450
		x"0A",x"34",x"63",x"66",x"BD",x"D8",x"79",x"DA", -- 0x3458
		x"E3",x"BF",x"28",x"00",x"18",x"74",x"62",x"28", -- 0x3460
		x"6A",x"8B",x"56",x"6A",x"50",x"1E",x"5D",x"73", -- 0x3468
		x"48",x"D5",x"87",x"44",x"53",x"18",x"7D",x"68", -- 0x3470
		x"C7",x"63",x"75",x"17",x"F3",x"05",x"4C",x"B4", -- 0x3478
		x"02",x"11",x"A4",x"27",x"F5",x"3B",x"2A",x"95", -- 0x3480
		x"B6",x"B5",x"F9",x"07",x"D5",x"7D",x"FE",x"19", -- 0x3488
		x"11",x"BF",x"7E",x"5D",x"4C",x"A3",x"B0",x"2D", -- 0x3490
		x"9F",x"E8",x"C8",x"F4",x"06",x"6C",x"F7",x"98", -- 0x3498
		x"8A",x"21",x"10",x"2C",x"9E",x"6D",x"DB",x"9A", -- 0x34A0
		x"E9",x"0A",x"28",x"02",x"64",x"CD",x"0E",x"26", -- 0x34A8
		x"AC",x"E5",x"A2",x"0B",x"8F",x"44",x"07",x"A4", -- 0x34B0
		x"D4",x"5C",x"9A",x"2C",x"B0",x"FE",x"96",x"8A", -- 0x34B8
		x"4E",x"8F",x"E4",x"A5",x"77",x"56",x"E7",x"CC", -- 0x34C0
		x"5F",x"83",x"7A",x"DB",x"3C",x"16",x"D3",x"23", -- 0x34C8
		x"7D",x"82",x"57",x"05",x"C9",x"80",x"CF",x"86", -- 0x34D0
		x"28",x"7C",x"EF",x"95",x"58",x"08",x"EF",x"A2", -- 0x34D8
		x"EB",x"A0",x"7F",x"18",x"B6",x"B8",x"6F",x"EC", -- 0x34E0
		x"2D",x"5B",x"C8",x"41",x"06",x"43",x"61",x"BF", -- 0x34E8
		x"8A",x"E3",x"92",x"C5",x"4F",x"5C",x"7C",x"B7", -- 0x34F0
		x"6F",x"EB",x"86",x"5D",x"5E",x"4A",x"6B",x"B8", -- 0x34F8
		x"96",x"73",x"BF",x"2F",x"57",x"72",x"CE",x"98", -- 0x3500
		x"A9",x"16",x"1D",x"1C",x"FF",x"18",x"8B",x"C7", -- 0x3508
		x"C9",x"C8",x"1A",x"66",x"FF",x"64",x"89",x"F9", -- 0x3510
		x"DB",x"D1",x"62",x"6C",x"64",x"C5",x"19",x"19", -- 0x3518
		x"8D",x"B4",x"C2",x"67",x"9D",x"20",x"DF",x"A6", -- 0x3520
		x"04",x"28",x"26",x"D9",x"2B",x"78",x"26",x"00", -- 0x3528
		x"3B",x"06",x"E7",x"B0",x"00",x"41",x"0F",x"63", -- 0x3530
		x"00",x"C0",x"4D",x"81",x"7C",x"D0",x"68",x"10", -- 0x3538
		x"04",x"E7",x"32",x"03",x"30",x"F8",x"3A",x"67", -- 0x3540
		x"4E",x"35",x"6C",x"7F",x"EB",x"87",x"6B",x"F7", -- 0x3548
		x"40",x"8A",x"BA",x"EB",x"E7",x"78",x"29",x"A4", -- 0x3550
		x"41",x"1A",x"BD",x"74",x"65",x"21",x"12",x"BC", -- 0x3558
		x"21",x"EB",x"CD",x"49",x"C1",x"FF",x"C4",x"14", -- 0x3560
		x"6E",x"32",x"71",x"26",x"F6",x"DE",x"C6",x"F2", -- 0x3568
		x"79",x"D0",x"E9",x"47",x"14",x"E0",x"C0",x"5C", -- 0x3570
		x"43",x"84",x"0B",x"DC",x"0C",x"B2",x"DE",x"EA", -- 0x3578
		x"AB",x"3C",x"40",x"3E",x"6C",x"99",x"ED",x"4F", -- 0x3580
		x"93",x"FB",x"60",x"0A",x"F5",x"0F",x"F5",x"B8", -- 0x3588
		x"11",x"69",x"1B",x"E8",x"2B",x"30",x"7D",x"63", -- 0x3590
		x"B0",x"D4",x"8C",x"17",x"18",x"8E",x"E6",x"43", -- 0x3598
		x"8B",x"48",x"33",x"9C",x"BA",x"3D",x"47",x"73", -- 0x35A0
		x"A5",x"04",x"0A",x"0F",x"1B",x"25",x"5D",x"15", -- 0x35A8
		x"FA",x"24",x"7C",x"13",x"03",x"2D",x"72",x"BE", -- 0x35B0
		x"64",x"5C",x"3F",x"F7",x"E4",x"59",x"09",x"79", -- 0x35B8
		x"0E",x"8C",x"7B",x"74",x"9D",x"9D",x"D5",x"4B", -- 0x35C0
		x"85",x"BB",x"5D",x"BF",x"4D",x"B9",x"A0",x"31", -- 0x35C8
		x"25",x"A5",x"D2",x"46",x"AF",x"09",x"DE",x"10", -- 0x35D0
		x"4B",x"CC",x"B3",x"67",x"94",x"CF",x"39",x"79", -- 0x35D8
		x"53",x"74",x"59",x"29",x"5A",x"5A",x"29",x"B4", -- 0x35E0
		x"4A",x"36",x"AB",x"48",x"C7",x"5F",x"13",x"80", -- 0x35E8
		x"B6",x"AA",x"D0",x"2C",x"28",x"C2",x"5E",x"53", -- 0x35F0
		x"88",x"1D",x"53",x"E1",x"DA",x"C8",x"E3",x"BC", -- 0x35F8
		x"34",x"E9",x"3D",x"FF",x"D1",x"A6",x"B6",x"BD", -- 0x3600
		x"CF",x"27",x"11",x"88",x"F9",x"55",x"0A",x"B9", -- 0x3608
		x"5F",x"0F",x"9D",x"11",x"E8",x"FF",x"E9",x"B3", -- 0x3610
		x"B3",x"14",x"06",x"C7",x"19",x"4D",x"CB",x"84", -- 0x3618
		x"17",x"A1",x"CF",x"B0",x"7F",x"65",x"AE",x"43", -- 0x3620
		x"6B",x"3B",x"41",x"AA",x"D7",x"E1",x"2F",x"E6", -- 0x3628
		x"20",x"64",x"6E",x"D7",x"F1",x"D3",x"19",x"37", -- 0x3630
		x"72",x"64",x"5F",x"49",x"43",x"0D",x"98",x"C0", -- 0x3638
		x"74",x"12",x"33",x"6E",x"76",x"AA",x"BC",x"E0", -- 0x3640
		x"D7",x"82",x"07",x"B8",x"F4",x"26",x"A6",x"B6", -- 0x3648
		x"8E",x"31",x"7D",x"50",x"D7",x"13",x"C7",x"77", -- 0x3650
		x"18",x"C6",x"3C",x"16",x"EE",x"BB",x"D2",x"ED", -- 0x3658
		x"97",x"2A",x"C7",x"9C",x"52",x"63",x"39",x"C0", -- 0x3660
		x"BA",x"7C",x"37",x"47",x"37",x"4D",x"99",x"25", -- 0x3668
		x"63",x"2A",x"BF",x"57",x"44",x"46",x"34",x"1E", -- 0x3670
		x"38",x"EC",x"19",x"B3",x"A9",x"CF",x"F3",x"0B", -- 0x3678
		x"6A",x"1C",x"DF",x"BF",x"16",x"38",x"4B",x"A3", -- 0x3680
		x"B0",x"BF",x"B0",x"E0",x"E4",x"29",x"61",x"E5", -- 0x3688
		x"AC",x"B6",x"C9",x"F0",x"6F",x"2F",x"C3",x"55", -- 0x3690
		x"B4",x"C9",x"CB",x"94",x"00",x"1A",x"BF",x"55", -- 0x3698
		x"72",x"5B",x"BD",x"2A",x"29",x"1A",x"BC",x"37", -- 0x36A0
		x"83",x"F6",x"BF",x"04",x"38",x"15",x"FE",x"2B", -- 0x36A8
		x"18",x"FA",x"85",x"04",x"B5",x"0D",x"69",x"61", -- 0x36B0
		x"06",x"38",x"CA",x"1F",x"8F",x"9C",x"D4",x"63", -- 0x36B8
		x"DB",x"74",x"EC",x"A9",x"E4",x"C4",x"15",x"01", -- 0x36C0
		x"67",x"89",x"73",x"8B",x"3D",x"BD",x"C3",x"A0", -- 0x36C8
		x"7E",x"89",x"DB",x"12",x"9F",x"01",x"36",x"02", -- 0x36D0
		x"CD",x"11",x"66",x"C7",x"AF",x"86",x"D5",x"91", -- 0x36D8
		x"E5",x"9E",x"F2",x"0E",x"C0",x"CD",x"48",x"F8", -- 0x36E0
		x"44",x"B2",x"0A",x"FC",x"1C",x"A1",x"7F",x"22", -- 0x36E8
		x"98",x"22",x"CC",x"0D",x"D7",x"26",x"44",x"18", -- 0x36F0
		x"75",x"83",x"33",x"50",x"D8",x"A1",x"BA",x"41", -- 0x36F8
		x"4D",x"47",x"26",x"80",x"E4",x"B0",x"7B",x"29", -- 0x3700
		x"F4",x"E0",x"9B",x"E2",x"AE",x"6B",x"99",x"E4", -- 0x3708
		x"11",x"C1",x"46",x"B5",x"FB",x"5D",x"BC",x"1D", -- 0x3710
		x"64",x"32",x"2D",x"4C",x"34",x"72",x"55",x"64", -- 0x3718
		x"63",x"08",x"A1",x"98",x"E4",x"AE",x"8B",x"BE", -- 0x3720
		x"70",x"70",x"AF",x"8F",x"75",x"DD",x"3D",x"29", -- 0x3728
		x"18",x"1A",x"22",x"BC",x"F7",x"35",x"C2",x"8B", -- 0x3730
		x"57",x"F0",x"2C",x"A0",x"3D",x"5B",x"84",x"AC", -- 0x3738
		x"85",x"96",x"7C",x"6F",x"5A",x"41",x"4D",x"AE", -- 0x3740
		x"15",x"6F",x"2E",x"E6",x"05",x"31",x"4C",x"DC", -- 0x3748
		x"FE",x"B3",x"3A",x"2E",x"C7",x"AE",x"B7",x"14", -- 0x3750
		x"5B",x"19",x"97",x"26",x"FE",x"ED",x"FB",x"4E", -- 0x3758
		x"4E",x"4D",x"3D",x"62",x"96",x"09",x"10",x"E9", -- 0x3760
		x"7C",x"AF",x"72",x"09",x"3C",x"C6",x"5C",x"CB", -- 0x3768
		x"7B",x"69",x"82",x"CB",x"47",x"4C",x"C0",x"35", -- 0x3770
		x"D7",x"39",x"28",x"7D",x"A0",x"F2",x"A6",x"B3", -- 0x3778
		x"3C",x"11",x"D3",x"FC",x"AD",x"42",x"A9",x"01", -- 0x3780
		x"B6",x"CC",x"9F",x"AE",x"B5",x"58",x"B2",x"DA", -- 0x3788
		x"54",x"CE",x"7C",x"81",x"FB",x"2D",x"3E",x"9A", -- 0x3790
		x"2F",x"80",x"B4",x"D5",x"48",x"59",x"90",x"3E", -- 0x3798
		x"BF",x"D7",x"9C",x"6A",x"E1",x"70",x"7B",x"F1", -- 0x37A0
		x"C2",x"56",x"E5",x"B7",x"29",x"2C",x"DE",x"2F", -- 0x37A8
		x"65",x"AC",x"CA",x"0F",x"D4",x"39",x"B8",x"B7", -- 0x37B0
		x"43",x"A2",x"1D",x"5F",x"42",x"C5",x"82",x"44", -- 0x37B8
		x"2F",x"A6",x"BC",x"48",x"51",x"F3",x"0C",x"11", -- 0x37C0
		x"CC",x"61",x"6D",x"B8",x"5A",x"46",x"7A",x"F6", -- 0x37C8
		x"BD",x"DF",x"66",x"92",x"82",x"AC",x"0F",x"95", -- 0x37D0
		x"42",x"D7",x"BE",x"0E",x"6F",x"65",x"17",x"08", -- 0x37D8
		x"D0",x"A2",x"A1",x"91",x"9B",x"EB",x"56",x"17", -- 0x37E0
		x"17",x"C4",x"2A",x"64",x"06",x"BF",x"1D",x"BE", -- 0x37E8
		x"42",x"41",x"41",x"EB",x"73",x"50",x"7F",x"AA", -- 0x37F0
		x"D4",x"23",x"CE",x"19",x"49",x"7B",x"23",x"20", -- 0x37F8
		x"ED",x"16",x"C2",x"7A",x"F8",x"16",x"72",x"D4", -- 0x3800
		x"07",x"95",x"CB",x"CC",x"91",x"A5",x"3F",x"58", -- 0x3808
		x"C5",x"FC",x"10",x"58",x"AA",x"7D",x"65",x"08", -- 0x3810
		x"ED",x"94",x"3D",x"59",x"FA",x"4C",x"A7",x"CF", -- 0x3818
		x"79",x"AF",x"FD",x"69",x"F3",x"D6",x"61",x"E1", -- 0x3820
		x"77",x"13",x"43",x"92",x"1F",x"0F",x"0C",x"7A", -- 0x3828
		x"AD",x"12",x"2F",x"7E",x"87",x"0E",x"CC",x"24", -- 0x3830
		x"88",x"C0",x"C3",x"D8",x"00",x"73",x"40",x"30", -- 0x3838
		x"FF",x"E3",x"5A",x"9D",x"19",x"17",x"76",x"02", -- 0x3840
		x"69",x"8F",x"B7",x"B2",x"26",x"96",x"2E",x"F4", -- 0x3848
		x"9E",x"01",x"DF",x"AA",x"7F",x"3E",x"B5",x"B7", -- 0x3850
		x"1E",x"A2",x"D9",x"52",x"E1",x"C9",x"8F",x"99", -- 0x3858
		x"01",x"05",x"5F",x"02",x"0B",x"47",x"6D",x"BD", -- 0x3860
		x"F7",x"83",x"9C",x"0E",x"47",x"CA",x"96",x"49", -- 0x3868
		x"B1",x"5F",x"8E",x"90",x"8D",x"98",x"77",x"63", -- 0x3870
		x"0C",x"1A",x"EF",x"42",x"BB",x"01",x"CB",x"3C", -- 0x3878
		x"EB",x"91",x"EB",x"54",x"57",x"B7",x"4D",x"30", -- 0x3880
		x"25",x"94",x"35",x"46",x"C1",x"2C",x"BB",x"AB", -- 0x3888
		x"AA",x"A7",x"A1",x"79",x"FB",x"A9",x"CC",x"74", -- 0x3890
		x"B0",x"18",x"7A",x"9F",x"E4",x"79",x"8C",x"14", -- 0x3898
		x"4C",x"AA",x"39",x"99",x"53",x"A6",x"AE",x"30", -- 0x38A0
		x"A4",x"73",x"4F",x"C7",x"71",x"8B",x"5C",x"8A", -- 0x38A8
		x"AD",x"C8",x"42",x"83",x"A2",x"5A",x"AD",x"04", -- 0x38B0
		x"0B",x"29",x"C8",x"11",x"18",x"C1",x"3E",x"AD", -- 0x38B8
		x"4E",x"CA",x"66",x"DD",x"DB",x"4A",x"EA",x"EE", -- 0x38C0
		x"AF",x"B6",x"D6",x"88",x"79",x"FC",x"EA",x"6B", -- 0x38C8
		x"87",x"90",x"71",x"18",x"BB",x"F0",x"17",x"47", -- 0x38D0
		x"FE",x"FA",x"F0",x"F5",x"0D",x"F9",x"09",x"7E", -- 0x38D8
		x"10",x"E9",x"E6",x"A7",x"C0",x"99",x"5C",x"E2", -- 0x38E0
		x"F9",x"C9",x"C6",x"90",x"40",x"91",x"CC",x"B5", -- 0x38E8
		x"20",x"6F",x"58",x"3B",x"D3",x"B5",x"73",x"23", -- 0x38F0
		x"96",x"92",x"84",x"B7",x"A8",x"65",x"81",x"7A", -- 0x38F8
		x"6F",x"BA",x"CF",x"B0",x"DB",x"26",x"EB",x"C0", -- 0x3900
		x"C5",x"54",x"DF",x"8D",x"B7",x"94",x"EF",x"4C", -- 0x3908
		x"0D",x"31",x"D2",x"6A",x"46",x"EF",x"31",x"E7", -- 0x3910
		x"2E",x"35",x"4B",x"E6",x"24",x"46",x"EF",x"30", -- 0x3918
		x"F5",x"0B",x"A8",x"74",x"40",x"5E",x"9D",x"AD", -- 0x3920
		x"90",x"57",x"4A",x"12",x"90",x"3C",x"04",x"E6", -- 0x3928
		x"3B",x"50",x"A4",x"54",x"CD",x"5F",x"3E",x"04", -- 0x3930
		x"64",x"60",x"B4",x"72",x"8D",x"C1",x"82",x"C6", -- 0x3938
		x"CB",x"96",x"AD",x"B2",x"DC",x"60",x"46",x"07", -- 0x3940
		x"47",x"E0",x"66",x"53",x"D8",x"AA",x"BD",x"EE", -- 0x3948
		x"42",x"57",x"81",x"A5",x"1F",x"11",x"93",x"B5", -- 0x3950
		x"35",x"4B",x"A0",x"57",x"E9",x"0F",x"30",x"4A", -- 0x3958
		x"40",x"D4",x"53",x"96",x"61",x"3F",x"99",x"B0", -- 0x3960
		x"A4",x"B1",x"59",x"B0",x"08",x"BE",x"13",x"D0", -- 0x3968
		x"9E",x"C1",x"09",x"65",x"1B",x"E1",x"75",x"9A", -- 0x3970
		x"C0",x"37",x"1C",x"FD",x"63",x"42",x"97",x"B7", -- 0x3978
		x"0F",x"30",x"63",x"65",x"41",x"3F",x"0A",x"20", -- 0x3980
		x"8E",x"21",x"9F",x"09",x"6B",x"88",x"99",x"50", -- 0x3988
		x"79",x"07",x"76",x"5F",x"F2",x"1D",x"95",x"41", -- 0x3990
		x"7A",x"FB",x"91",x"5F",x"E0",x"F0",x"D8",x"71", -- 0x3998
		x"B5",x"6D",x"39",x"0C",x"26",x"FB",x"06",x"D9", -- 0x39A0
		x"95",x"C9",x"E8",x"DD",x"EB",x"F1",x"1E",x"41", -- 0x39A8
		x"45",x"06",x"8B",x"93",x"0C",x"4C",x"90",x"F3", -- 0x39B0
		x"E4",x"E4",x"C3",x"23",x"16",x"00",x"09",x"A8", -- 0x39B8
		x"51",x"3B",x"F3",x"7E",x"E5",x"E9",x"6C",x"A4", -- 0x39C0
		x"70",x"01",x"AE",x"68",x"E0",x"98",x"BF",x"9F", -- 0x39C8
		x"85",x"5E",x"97",x"ED",x"3A",x"52",x"F0",x"90", -- 0x39D0
		x"C5",x"66",x"BB",x"F3",x"F9",x"E1",x"C6",x"EB", -- 0x39D8
		x"AE",x"D2",x"57",x"40",x"2A",x"01",x"0E",x"DE", -- 0x39E0
		x"14",x"8D",x"79",x"1E",x"A3",x"E2",x"B1",x"94", -- 0x39E8
		x"3C",x"96",x"84",x"AC",x"B3",x"93",x"54",x"7D", -- 0x39F0
		x"65",x"91",x"08",x"AB",x"40",x"D2",x"40",x"88", -- 0x39F8
		x"06",x"4D",x"5C",x"C0",x"96",x"D8",x"DB",x"87", -- 0x3A00
		x"7D",x"9A",x"55",x"39",x"E7",x"DA",x"CF",x"F1", -- 0x3A08
		x"53",x"65",x"EF",x"31",x"EF",x"50",x"B0",x"A1", -- 0x3A10
		x"F9",x"59",x"B7",x"1B",x"5F",x"D4",x"FC",x"D9", -- 0x3A18
		x"8A",x"F7",x"8F",x"B3",x"4D",x"40",x"AB",x"18", -- 0x3A20
		x"F9",x"57",x"49",x"01",x"3D",x"1A",x"83",x"56", -- 0x3A28
		x"A5",x"95",x"54",x"05",x"31",x"66",x"B5",x"A8", -- 0x3A30
		x"98",x"A4",x"77",x"4C",x"91",x"94",x"90",x"C9", -- 0x3A38
		x"16",x"E9",x"DA",x"18",x"DB",x"55",x"FA",x"FE", -- 0x3A40
		x"16",x"29",x"9F",x"82",x"D9",x"AC",x"E3",x"26", -- 0x3A48
		x"77",x"16",x"18",x"49",x"08",x"17",x"BF",x"BD", -- 0x3A50
		x"9B",x"9F",x"69",x"1E",x"CE",x"89",x"37",x"98", -- 0x3A58
		x"D1",x"8F",x"7C",x"C1",x"C4",x"D4",x"2D",x"74", -- 0x3A60
		x"6A",x"31",x"D0",x"71",x"F0",x"D1",x"78",x"12", -- 0x3A68
		x"54",x"64",x"35",x"09",x"A1",x"A3",x"65",x"57", -- 0x3A70
		x"E5",x"4C",x"17",x"76",x"18",x"CD",x"22",x"85", -- 0x3A78
		x"5F",x"05",x"0B",x"B1",x"15",x"20",x"87",x"9C", -- 0x3A80
		x"FD",x"68",x"B8",x"96",x"7E",x"DE",x"52",x"ED", -- 0x3A88
		x"49",x"1B",x"77",x"B9",x"7A",x"55",x"20",x"58", -- 0x3A90
		x"2F",x"EB",x"68",x"56",x"71",x"9A",x"5B",x"3A", -- 0x3A98
		x"97",x"08",x"84",x"D5",x"EB",x"F9",x"CF",x"56", -- 0x3AA0
		x"EF",x"43",x"76",x"F4",x"D3",x"9C",x"47",x"67", -- 0x3AA8
		x"29",x"9D",x"A2",x"55",x"B8",x"3C",x"CC",x"8D", -- 0x3AB0
		x"8D",x"B5",x"B0",x"44",x"E4",x"83",x"05",x"A9", -- 0x3AB8
		x"F1",x"CF",x"7D",x"A3",x"24",x"32",x"D1",x"09", -- 0x3AC0
		x"2E",x"4D",x"5F",x"86",x"8B",x"71",x"14",x"1B", -- 0x3AC8
		x"48",x"91",x"F6",x"21",x"BD",x"27",x"EB",x"8D", -- 0x3AD0
		x"11",x"A3",x"5A",x"FD",x"6F",x"73",x"04",x"63", -- 0x3AD8
		x"F4",x"B3",x"5C",x"5A",x"F7",x"0D",x"B8",x"7F", -- 0x3AE0
		x"C7",x"53",x"FB",x"EB",x"9B",x"14",x"90",x"F7", -- 0x3AE8
		x"89",x"E6",x"76",x"A8",x"43",x"12",x"DF",x"8A", -- 0x3AF0
		x"08",x"2A",x"E1",x"34",x"51",x"12",x"FB",x"1D", -- 0x3AF8
		x"A5",x"6C",x"A5",x"5A",x"2F",x"C4",x"CE",x"CA", -- 0x3B00
		x"46",x"67",x"0A",x"5D",x"17",x"3D",x"A1",x"0D", -- 0x3B08
		x"18",x"1F",x"5D",x"CC",x"89",x"11",x"D6",x"AF", -- 0x3B10
		x"93",x"94",x"E3",x"49",x"FB",x"9A",x"88",x"40", -- 0x3B18
		x"07",x"E2",x"08",x"7D",x"56",x"94",x"87",x"B7", -- 0x3B20
		x"62",x"9B",x"65",x"40",x"B8",x"71",x"A0",x"46", -- 0x3B28
		x"18",x"34",x"AA",x"E1",x"13",x"1D",x"86",x"55", -- 0x3B30
		x"F1",x"53",x"73",x"49",x"E5",x"00",x"1A",x"A6", -- 0x3B38
		x"EA",x"42",x"D2",x"60",x"74",x"DC",x"DB",x"99", -- 0x3B40
		x"A2",x"4B",x"79",x"E2",x"DA",x"B2",x"A5",x"E3", -- 0x3B48
		x"0A",x"72",x"78",x"BE",x"61",x"9A",x"7E",x"61", -- 0x3B50
		x"87",x"77",x"E9",x"AB",x"5D",x"BE",x"73",x"74", -- 0x3B58
		x"AE",x"A2",x"D7",x"B1",x"36",x"97",x"C9",x"A8", -- 0x3B60
		x"D6",x"99",x"0F",x"A0",x"19",x"82",x"00",x"10", -- 0x3B68
		x"D8",x"9A",x"50",x"F5",x"71",x"20",x"1E",x"5E", -- 0x3B70
		x"E4",x"32",x"3C",x"35",x"51",x"C9",x"4C",x"9F", -- 0x3B78
		x"9B",x"19",x"FB",x"41",x"05",x"CA",x"DE",x"8A", -- 0x3B80
		x"7B",x"09",x"27",x"74",x"C2",x"09",x"D4",x"69", -- 0x3B88
		x"30",x"D6",x"A1",x"A9",x"F8",x"87",x"4F",x"7A", -- 0x3B90
		x"95",x"4C",x"8A",x"E7",x"EB",x"62",x"FF",x"B7", -- 0x3B98
		x"48",x"6C",x"EC",x"6A",x"1B",x"95",x"A2",x"6C", -- 0x3BA0
		x"E6",x"CA",x"02",x"3B",x"A8",x"44",x"50",x"EE", -- 0x3BA8
		x"04",x"E0",x"0E",x"55",x"B4",x"D8",x"1F",x"3E", -- 0x3BB0
		x"91",x"86",x"5C",x"3D",x"C0",x"65",x"96",x"32", -- 0x3BB8
		x"4D",x"ED",x"B6",x"6D",x"98",x"3E",x"73",x"F1", -- 0x3BC0
		x"61",x"D6",x"15",x"17",x"27",x"B4",x"2A",x"4F", -- 0x3BC8
		x"F2",x"3E",x"0E",x"6C",x"65",x"E9",x"A5",x"01", -- 0x3BD0
		x"74",x"9F",x"E1",x"23",x"7B",x"59",x"E9",x"98", -- 0x3BD8
		x"8F",x"C4",x"2B",x"C7",x"66",x"CF",x"CE",x"46", -- 0x3BE0
		x"D4",x"99",x"86",x"44",x"30",x"F9",x"6C",x"C1", -- 0x3BE8
		x"6C",x"C4",x"87",x"A3",x"C7",x"85",x"E1",x"9C", -- 0x3BF0
		x"2B",x"80",x"D5",x"1C",x"09",x"67",x"2A",x"08", -- 0x3BF8
		x"75",x"9A",x"DB",x"A6",x"D6",x"B3",x"CE",x"0B", -- 0x3C00
		x"FD",x"7A",x"E0",x"90",x"C2",x"41",x"BF",x"8F", -- 0x3C08
		x"A6",x"C6",x"95",x"14",x"0C",x"B7",x"73",x"E2", -- 0x3C10
		x"EE",x"34",x"BE",x"5E",x"2A",x"88",x"82",x"45", -- 0x3C18
		x"70",x"98",x"21",x"A8",x"7B",x"55",x"2C",x"3E", -- 0x3C20
		x"18",x"96",x"92",x"18",x"28",x"8A",x"E8",x"60", -- 0x3C28
		x"09",x"DC",x"FE",x"90",x"8E",x"2E",x"8E",x"00", -- 0x3C30
		x"17",x"34",x"2C",x"7E",x"10",x"61",x"1D",x"03", -- 0x3C38
		x"4F",x"45",x"DB",x"09",x"CD",x"4A",x"AB",x"AF", -- 0x3C40
		x"82",x"92",x"4A",x"6D",x"DF",x"BA",x"7E",x"C6", -- 0x3C48
		x"57",x"4A",x"E8",x"0D",x"15",x"E8",x"E5",x"D1", -- 0x3C50
		x"F1",x"FC",x"C8",x"5F",x"33",x"C7",x"3C",x"B0", -- 0x3C58
		x"67",x"BD",x"2C",x"CF",x"A9",x"E0",x"7C",x"B4", -- 0x3C60
		x"4F",x"F1",x"55",x"80",x"F1",x"5B",x"A2",x"C6", -- 0x3C68
		x"16",x"74",x"A8",x"F4",x"49",x"DE",x"50",x"A1", -- 0x3C70
		x"28",x"64",x"B3",x"28",x"2D",x"0B",x"D0",x"C3", -- 0x3C78
		x"DB",x"63",x"FF",x"63",x"B4",x"35",x"C3",x"6B", -- 0x3C80
		x"FE",x"5B",x"34",x"4F",x"E1",x"16",x"71",x"CA", -- 0x3C88
		x"D0",x"30",x"D6",x"38",x"6F",x"6E",x"6B",x"CD", -- 0x3C90
		x"DC",x"AE",x"8D",x"F4",x"9F",x"32",x"3F",x"14", -- 0x3C98
		x"3A",x"F9",x"45",x"76",x"80",x"C4",x"52",x"AF", -- 0x3CA0
		x"AC",x"C9",x"0F",x"0D",x"0D",x"67",x"08",x"E0", -- 0x3CA8
		x"AF",x"A6",x"85",x"02",x"87",x"7C",x"4A",x"8C", -- 0x3CB0
		x"86",x"A2",x"AB",x"A0",x"89",x"00",x"3B",x"C4", -- 0x3CB8
		x"53",x"D1",x"9B",x"A1",x"1D",x"88",x"EB",x"CD", -- 0x3CC0
		x"BD",x"28",x"4D",x"DA",x"7B",x"0D",x"1E",x"4E", -- 0x3CC8
		x"58",x"99",x"FC",x"C2",x"4F",x"E9",x"B7",x"3A", -- 0x3CD0
		x"B9",x"F8",x"73",x"FC",x"3E",x"B7",x"59",x"96", -- 0x3CD8
		x"42",x"3B",x"47",x"99",x"7F",x"10",x"1B",x"51", -- 0x3CE0
		x"09",x"D9",x"E2",x"15",x"99",x"CC",x"5B",x"DB", -- 0x3CE8
		x"F1",x"01",x"11",x"A5",x"02",x"10",x"F7",x"79", -- 0x3CF0
		x"29",x"14",x"01",x"09",x"6F",x"E6",x"EC",x"BB", -- 0x3CF8
		x"CA",x"F5",x"2B",x"CE",x"2A",x"66",x"FD",x"2B", -- 0x3D00
		x"BB",x"5C",x"50",x"96",x"3A",x"A6",x"67",x"F2", -- 0x3D08
		x"A5",x"ED",x"F7",x"5B",x"4E",x"D4",x"E8",x"02", -- 0x3D10
		x"77",x"50",x"B9",x"A1",x"78",x"83",x"42",x"95", -- 0x3D18
		x"EA",x"99",x"C9",x"2B",x"8B",x"BA",x"28",x"8C", -- 0x3D20
		x"59",x"07",x"0D",x"1D",x"66",x"D1",x"E4",x"CE", -- 0x3D28
		x"01",x"C7",x"4A",x"B0",x"4F",x"66",x"5A",x"CC", -- 0x3D30
		x"81",x"22",x"83",x"B5",x"4C",x"C6",x"DF",x"2D", -- 0x3D38
		x"81",x"17",x"6A",x"A2",x"DD",x"E5",x"ED",x"51", -- 0x3D40
		x"59",x"8A",x"F9",x"03",x"F5",x"8D",x"1A",x"CB", -- 0x3D48
		x"91",x"D3",x"AD",x"3F",x"7C",x"BD",x"AF",x"12", -- 0x3D50
		x"51",x"00",x"39",x"08",x"E5",x"AD",x"92",x"49", -- 0x3D58
		x"07",x"21",x"8D",x"D5",x"74",x"AD",x"93",x"7A", -- 0x3D60
		x"21",x"8C",x"50",x"72",x"7E",x"D5",x"00",x"E9", -- 0x3D68
		x"48",x"A1",x"99",x"4A",x"A0",x"30",x"97",x"C8", -- 0x3D70
		x"C6",x"70",x"6F",x"0E",x"68",x"73",x"AD",x"FC", -- 0x3D78
		x"A4",x"CC",x"5B",x"FA",x"B2",x"72",x"F9",x"D4", -- 0x3D80
		x"5B",x"B2",x"BF",x"C9",x"82",x"19",x"0E",x"CA", -- 0x3D88
		x"DF",x"D1",x"FB",x"18",x"7F",x"11",x"F6",x"B9", -- 0x3D90
		x"7B",x"8E",x"E1",x"4E",x"B8",x"08",x"77",x"D0", -- 0x3D98
		x"5E",x"5A",x"BF",x"C2",x"4F",x"59",x"A5",x"18", -- 0x3DA0
		x"A4",x"EB",x"DF",x"55",x"49",x"6E",x"F1",x"78", -- 0x3DA8
		x"45",x"85",x"BD",x"41",x"C6",x"CA",x"71",x"53", -- 0x3DB0
		x"33",x"04",x"1F",x"33",x"70",x"EF",x"5A",x"A8", -- 0x3DB8
		x"7C",x"2A",x"37",x"4F",x"83",x"CB",x"AF",x"C5", -- 0x3DC0
		x"A9",x"F3",x"E2",x"60",x"3B",x"EA",x"EB",x"C1", -- 0x3DC8
		x"7B",x"D6",x"F9",x"9A",x"3B",x"07",x"5C",x"9E", -- 0x3DD0
		x"17",x"16",x"F5",x"9E",x"DD",x"6E",x"12",x"9C", -- 0x3DD8
		x"37",x"4E",x"DB",x"CA",x"7A",x"9A",x"A2",x"DC", -- 0x3DE0
		x"63",x"C4",x"34",x"0D",x"41",x"FE",x"BD",x"AD", -- 0x3DE8
		x"C9",x"6F",x"76",x"F4",x"AD",x"15",x"CB",x"49", -- 0x3DF0
		x"B4",x"27",x"33",x"52",x"E0",x"87",x"99",x"9A", -- 0x3DF8
		x"3F",x"F9",x"D7",x"CA",x"7C",x"97",x"51",x"15", -- 0x3E00
		x"78",x"1D",x"DE",x"5B",x"2F",x"DE",x"96",x"DC", -- 0x3E08
		x"8E",x"6B",x"B9",x"3E",x"DA",x"77",x"FB",x"46", -- 0x3E10
		x"37",x"A6",x"88",x"74",x"C1",x"D5",x"C3",x"F2", -- 0x3E18
		x"C5",x"1C",x"EA",x"27",x"DC",x"35",x"12",x"9C", -- 0x3E20
		x"D1",x"BD",x"7E",x"08",x"43",x"BF",x"45",x"B4", -- 0x3E28
		x"E6",x"F1",x"78",x"6D",x"2B",x"CE",x"B6",x"D2", -- 0x3E30
		x"26",x"7B",x"6A",x"69",x"D5",x"01",x"A7",x"18", -- 0x3E38
		x"76",x"15",x"99",x"6F",x"5F",x"55",x"7B",x"D3", -- 0x3E40
		x"21",x"63",x"08",x"F7",x"F1",x"28",x"19",x"F4", -- 0x3E48
		x"D1",x"02",x"C5",x"A4",x"D2",x"46",x"E0",x"62", -- 0x3E50
		x"75",x"2E",x"E4",x"F7",x"42",x"26",x"A7",x"73", -- 0x3E58
		x"6A",x"0E",x"44",x"3C",x"36",x"66",x"58",x"A4", -- 0x3E60
		x"2C",x"B2",x"41",x"9B",x"37",x"3C",x"D5",x"D4", -- 0x3E68
		x"48",x"3D",x"C0",x"4E",x"38",x"DC",x"E7",x"16", -- 0x3E70
		x"6B",x"8E",x"61",x"15",x"20",x"6B",x"D9",x"40", -- 0x3E78
		x"C7",x"2E",x"E3",x"3D",x"7F",x"E9",x"55",x"6C", -- 0x3E80
		x"33",x"64",x"FE",x"87",x"CD",x"C8",x"57",x"49", -- 0x3E88
		x"4B",x"CA",x"83",x"9D",x"13",x"64",x"C7",x"25", -- 0x3E90
		x"BE",x"9A",x"2F",x"F7",x"36",x"0E",x"DA",x"43", -- 0x3E98
		x"CC",x"44",x"84",x"A0",x"14",x"E1",x"23",x"4D", -- 0x3EA0
		x"AD",x"31",x"CA",x"4F",x"2E",x"00",x"D7",x"22", -- 0x3EA8
		x"B8",x"05",x"E3",x"18",x"64",x"19",x"24",x"04", -- 0x3EB0
		x"59",x"5A",x"72",x"21",x"86",x"57",x"41",x"C5", -- 0x3EB8
		x"4F",x"69",x"87",x"CE",x"FB",x"3D",x"E1",x"3D", -- 0x3EC0
		x"25",x"D7",x"6B",x"B9",x"A0",x"50",x"C3",x"31", -- 0x3EC8
		x"02",x"13",x"C3",x"A3",x"C4",x"29",x"1D",x"FD", -- 0x3ED0
		x"DF",x"59",x"3C",x"F7",x"1F",x"59",x"BB",x"FA", -- 0x3ED8
		x"96",x"E5",x"AB",x"C7",x"69",x"14",x"3A",x"FB", -- 0x3EE0
		x"D2",x"91",x"4B",x"F1",x"76",x"78",x"A7",x"9F", -- 0x3EE8
		x"BB",x"D5",x"57",x"32",x"A4",x"62",x"D6",x"9F", -- 0x3EF0
		x"03",x"B4",x"70",x"B1",x"9A",x"B4",x"4A",x"12", -- 0x3EF8
		x"55",x"10",x"C1",x"67",x"2B",x"2F",x"31",x"DF", -- 0x3F00
		x"F0",x"58",x"AB",x"A6",x"D3",x"98",x"F6",x"D6", -- 0x3F08
		x"52",x"47",x"E8",x"4D",x"63",x"BA",x"F6",x"B4", -- 0x3F10
		x"B6",x"43",x"74",x"28",x"C7",x"A9",x"23",x"FD", -- 0x3F18
		x"F8",x"3B",x"88",x"68",x"20",x"EA",x"53",x"A0", -- 0x3F20
		x"8B",x"11",x"ED",x"7C",x"16",x"36",x"29",x"DD", -- 0x3F28
		x"5A",x"70",x"08",x"DF",x"2C",x"54",x"78",x"15", -- 0x3F30
		x"1D",x"D4",x"07",x"12",x"01",x"BB",x"2A",x"9D", -- 0x3F38
		x"CF",x"DB",x"49",x"B7",x"43",x"01",x"93",x"8D", -- 0x3F40
		x"10",x"87",x"1B",x"A1",x"E8",x"33",x"FB",x"75", -- 0x3F48
		x"F8",x"3B",x"C2",x"E1",x"34",x"FE",x"5E",x"9D", -- 0x3F50
		x"A8",x"38",x"2A",x"25",x"32",x"A6",x"9D",x"C6", -- 0x3F58
		x"49",x"43",x"79",x"37",x"F3",x"6D",x"B4",x"71", -- 0x3F60
		x"AE",x"50",x"92",x"63",x"D1",x"24",x"12",x"CF", -- 0x3F68
		x"54",x"26",x"D9",x"8B",x"8A",x"D0",x"B5",x"02", -- 0x3F70
		x"B4",x"00",x"A9",x"F9",x"A5",x"65",x"83",x"64", -- 0x3F78
		x"EB",x"1C",x"6B",x"33",x"7C",x"13",x"15",x"5D", -- 0x3F80
		x"E4",x"06",x"C9",x"81",x"94",x"93",x"F2",x"E7", -- 0x3F88
		x"8D",x"1B",x"E4",x"CF",x"DE",x"0E",x"5F",x"24", -- 0x3F90
		x"B5",x"F1",x"27",x"62",x"7A",x"9E",x"7C",x"D1", -- 0x3F98
		x"3C",x"8E",x"F2",x"57",x"8F",x"CB",x"7B",x"C6", -- 0x3FA0
		x"B3",x"20",x"04",x"A3",x"B2",x"0B",x"7D",x"28", -- 0x3FA8
		x"9F",x"8C",x"31",x"F9",x"DA",x"D4",x"82",x"58", -- 0x3FB0
		x"DB",x"16",x"27",x"31",x"98",x"38",x"2F",x"55", -- 0x3FB8
		x"68",x"E0",x"14",x"D3",x"01",x"AD",x"32",x"F0", -- 0x3FC0
		x"8A",x"31",x"F7",x"AE",x"45",x"ED",x"2A",x"FC", -- 0x3FC8
		x"E9",x"C6",x"8E",x"42",x"96",x"DF",x"57",x"26", -- 0x3FD0
		x"38",x"D0",x"9F",x"2C",x"A1",x"65",x"7D",x"49", -- 0x3FD8
		x"B1",x"18",x"97",x"EC",x"94",x"4A",x"B5",x"2F", -- 0x3FE0
		x"F3",x"2F",x"D4",x"39",x"CE",x"69",x"42",x"0E", -- 0x3FE8
		x"71",x"88",x"DB",x"A5",x"DC",x"BD",x"C5",x"FB", -- 0x3FF0
		x"25",x"75",x"22",x"61",x"33",x"95",x"F4",x"81"  -- 0x3FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
