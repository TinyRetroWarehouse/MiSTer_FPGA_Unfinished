-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_A1 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_A1 is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"04",x"00",x"10",x"3C",x"1E",x"0E",x"04",x"05", -- 0x0000
		x"81",x"80",x"50",x"B8",x"FC",x"DD",x"CE",x"EE", -- 0x0008
		x"00",x"04",x"00",x"00",x"08",x"0C",x"0E",x"06", -- 0x0010
		x"82",x"00",x"00",x"00",x"60",x"DC",x"CE",x"67", -- 0x0018
		x"81",x"C0",x"40",x"80",x"B0",x"99",x"DB",x"B1", -- 0x0020
		x"F8",x"B8",x"56",x"46",x"62",x"81",x"83",x"4F", -- 0x0028
		x"00",x"00",x"00",x"08",x"00",x"80",x"C2",x"C0", -- 0x0030
		x"E1",x"47",x"8C",x"C2",x"45",x"CF",x"A9",x"F3", -- 0x0038
		x"00",x"80",x"60",x"F0",x"F0",x"A0",x"B3",x"87", -- 0x0040
		x"C7",x"C3",x"E3",x"48",x"F8",x"E2",x"77",x"BF", -- 0x0048
		x"00",x"C0",x"E0",x"40",x"00",x"00",x"00",x"80", -- 0x0050
		x"80",x"30",x"78",x"38",x"18",x"04",x"08",x"CF", -- 0x0058
		x"80",x"00",x"60",x"60",x"F0",x"60",x"40",x"9C", -- 0x0060
		x"9C",x"BE",x"6E",x"34",x"10",x"1E",x"BE",x"EF", -- 0x0068
		x"00",x"00",x"00",x"10",x"38",x"28",x"18",x"00", -- 0x0070
		x"02",x"00",x"00",x"30",x"38",x"18",x"00",x"00", -- 0x0078
		x"00",x"40",x"00",x"18",x"0C",x"1C",x"1C",x"00", -- 0x0080
		x"80",x"80",x"4C",x"5C",x"6E",x"96",x"8F",x"4F", -- 0x0088
		x"00",x"00",x"10",x"00",x"00",x"04",x"06",x"06", -- 0x0090
		x"30",x"78",x"1C",x"3C",x"18",x"18",x"00",x"00", -- 0x0098
		x"DF",x"B7",x"32",x"70",x"BA",x"57",x"E7",x"E6", -- 0x00A0
		x"EA",x"87",x"43",x"E2",x"E1",x"F5",x"DE",x"EE", -- 0x00A8
		x"00",x"0C",x"1E",x"06",x"8E",x"C7",x"42",x"80", -- 0x00B0
		x"80",x"04",x"40",x"E0",x"40",x"D4",x"CE",x"E6", -- 0x00B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x00C0
		x"00",x"00",x"00",x"04",x"0F",x"27",x"1E",x"EE", -- 0x00C8
		x"00",x"00",x"00",x"00",x"40",x"E0",x"E0",x"40", -- 0x00D0
		x"21",x"03",x"07",x"03",x"62",x"D5",x"DF",x"E7", -- 0x00D8
		x"00",x"40",x"00",x"00",x"03",x"07",x"07",x"0F", -- 0x00E0
		x"DB",x"CB",x"E1",x"40",x"F0",x"E0",x"74",x"BE", -- 0x00E8
		x"01",x"07",x"07",x"19",x"1E",x"3F",x"8F",x"9F", -- 0x00F0
		x"CA",x"5D",x"17",x"0F",x"1B",x"06",x"09",x"CF", -- 0x00F8
		x"10",x"30",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0100
		x"03",x"00",x"01",x"08",x"18",x"2E",x"3F",x"0F", -- 0x0108
		x"01",x"01",x"03",x"09",x"1E",x"07",x"0F",x"85", -- 0x0110
		x"80",x"C1",x"8B",x"1F",x"0F",x"76",x"09",x"CF", -- 0x0118
		x"00",x"01",x"01",x"03",x"00",x"00",x"00",x"18", -- 0x0120
		x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0128
		x"01",x"83",x"CD",x"CD",x"8E",x"07",x"05",x"0A", -- 0x0130
		x"1A",x"39",x"14",x"0A",x"2D",x"77",x"79",x"BB", -- 0x0138
		x"00",x"20",x"00",x"00",x"08",x"3C",x"1C",x"0E", -- 0x0140
		x"1E",x"0C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0148
		x"00",x"06",x"03",x"10",x"28",x"18",x"00",x"00", -- 0x0150
		x"02",x"01",x"00",x"0A",x"1D",x"1F",x"09",x"1B", -- 0x0158
		x"00",x"30",x"00",x"00",x"00",x"00",x"05",x"07", -- 0x0160
		x"0E",x"07",x"0B",x"02",x"20",x"60",x"7E",x"2E", -- 0x0168
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"15",x"0B", -- 0x0170
		x"87",x"A7",x"B7",x"53",x"62",x"D5",x"DF",x"E7", -- 0x0178
		x"9F",x"C3",x"45",x"8F",x"87",x"8B",x"44",x"20", -- 0x0180
		x"00",x"03",x"03",x"03",x"01",x"00",x"00",x"00", -- 0x0188
		x"CE",x"B2",x"10",x"80",x"00",x"00",x"18",x"1C", -- 0x0190
		x"1C",x"08",x"00",x"80",x"80",x"80",x"00",x"00", -- 0x0198
		x"1F",x"8F",x"6C",x"F1",x"F8",x"A9",x"B1",x"98", -- 0x01A0
		x"D8",x"F0",x"F8",x"50",x"E0",x"60",x"00",x"00", -- 0x01A8
		x"EF",x"AB",x"C3",x"61",x"60",x"21",x"89",x"9C", -- 0x01B0
		x"88",x"1C",x"1C",x"08",x"00",x"00",x"00",x"00", -- 0x01B8
		x"2E",x"47",x"17",x"1C",x"DD",x"79",x"79",x"38", -- 0x01C0
		x"90",x"F8",x"68",x"30",x"70",x"60",x"00",x"00", -- 0x01C8
		x"19",x"3E",x"3E",x"94",x"84",x"80",x"60",x"E0", -- 0x01D0
		x"40",x"18",x"1C",x"1C",x"1C",x"0C",x"08",x"00", -- 0x01D8
		x"EF",x"47",x"02",x"00",x"C0",x"70",x"78",x"B8", -- 0x01E0
		x"90",x"D8",x"60",x"30",x"70",x"20",x"80",x"80", -- 0x01E8
		x"00",x"00",x"10",x"08",x"18",x"1C",x"08",x"00", -- 0x01F0
		x"00",x"00",x"30",x"78",x"38",x"18",x"00",x"00", -- 0x01F8
		x"EE",x"46",x"06",x"40",x"E0",x"70",x"20",x"00", -- 0x0200
		x"0C",x"0E",x"06",x"00",x"00",x"00",x"00",x"00", -- 0x0208
		x"00",x"00",x"30",x"78",x"38",x"58",x"00",x"00", -- 0x0210
		x"00",x"00",x"02",x"03",x"C0",x"60",x"00",x"00", -- 0x0218
		x"1F",x"97",x"72",x"F2",x"F0",x"B8",x"B0",x"91", -- 0x0220
		x"D3",x"C3",x"E7",x"4D",x"E5",x"E0",x"70",x"BE", -- 0x0228
		x"C4",x"80",x"10",x"18",x"38",x"18",x"00",x"80", -- 0x0230
		x"C0",x"40",x"E0",x"C0",x"00",x"02",x"02",x"00", -- 0x0238
		x"3F",x"1F",x"0D",x"03",x"06",x"00",x"00",x"00", -- 0x0240
		x"00",x"02",x"07",x"07",x"02",x"00",x"00",x"00", -- 0x0248
		x"F7",x"AB",x"D3",x"E1",x"52",x"05",x"0F",x"06", -- 0x0250
		x"02",x"00",x"00",x"80",x"00",x"00",x"00",x"00", -- 0x0258
		x"EE",x"47",x"05",x"00",x"C0",x"70",x"79",x"3B", -- 0x0260
		x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0268
		x"19",x"BE",x"FF",x"DF",x"17",x"06",x"C4",x"D0", -- 0x0270
		x"5C",x"06",x"0E",x"03",x"C3",x"65",x"C0",x"00", -- 0x0278
		x"4F",x"26",x"07",x"00",x"00",x"10",x"28",x"18", -- 0x0280
		x"1A",x"0E",x"0C",x"1C",x"0C",x"00",x"00",x"00", -- 0x0288
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"D5",x"6B", -- 0x0290
		x"FF",x"57",x"27",x"03",x"02",x"01",x"00",x"00", -- 0x0298
		x"00",x"00",x"00",x"01",x"01",x"03",x"01",x"00", -- 0x02A0
		x"03",x"03",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x02A8
		x"17",x"0B",x"53",x"21",x"22",x"C1",x"B7",x"C1", -- 0x02B0
		x"C0",x"01",x"C1",x"C1",x"80",x"00",x"00",x"00", -- 0x02B8
		x"00",x"60",x"60",x"00",x"04",x"06",x"06",x"00", -- 0x02C0
		x"00",x"00",x"01",x"01",x"00",x"20",x"00",x"00", -- 0x02C8
		x"49",x"33",x"05",x"01",x"02",x"03",x"01",x"60", -- 0x02D0
		x"F0",x"B8",x"DC",x"8C",x"80",x"00",x"00",x"00", -- 0x02D8
		x"5F",x"3E",x"34",x"00",x"0C",x"0E",x"07",x"07", -- 0x02E0
		x"0F",x"05",x"03",x"02",x"00",x"00",x"00",x"00", -- 0x02E8
		x"5F",x"67",x"2B",x"3F",x"5F",x"15",x"01",x"0B", -- 0x02F0
		x"9F",x"97",x"87",x"23",x"3A",x"5D",x"5F",x"27", -- 0x02F8
		x"00",x"20",x"31",x"00",x"03",x"00",x"00",x"00", -- 0x0300
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0308
		x"5F",x"E7",x"EB",x"DF",x"CF",x"C5",x"05",x"0B", -- 0x0310
		x"1F",x"77",x"77",x"93",x"62",x"75",x"5F",x"27", -- 0x0318
		x"DF",x"BF",x"35",x"74",x"B8",x"56",x"EC",x"F6", -- 0x0320
		x"C4",x"80",x"42",x"E2",x"F1",x"E1",x"DC",x"EC", -- 0x0328
		x"00",x"80",x"00",x"00",x"40",x"E1",x"62",x"C0", -- 0x0330
		x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0338
		x"EE",x"4F",x"13",x"10",x"C1",x"71",x"31",x"06", -- 0x0340
		x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0348
		x"19",x"3E",x"3F",x"DF",x"D7",x"EA",x"C0",x"C0", -- 0x0350
		x"80",x"00",x"00",x"40",x"C0",x"00",x"00",x"00", -- 0x0358
		x"20",x"30",x"00",x"00",x"00",x"08",x"0C",x"06", -- 0x0360
		x"8E",x"C6",x"E4",x"E0",x"63",x"73",x"BA",x"ED", -- 0x0368
		x"00",x"00",x"00",x"00",x"20",x"30",x"F0",x"7A", -- 0x0370
		x"5B",x"33",x"02",x"41",x"13",x"B9",x"74",x"7E", -- 0x0378
		x"00",x"01",x"09",x"1E",x"0C",x"1C",x"0B",x"07", -- 0x0380
		x"0B",x"01",x"00",x"0C",x"0A",x"06",x"00",x"00", -- 0x0388
		x"00",x"80",x"00",x"06",x"03",x"00",x"00",x"80", -- 0x0390
		x"80",x"00",x"00",x"2C",x"14",x"0E",x"04",x"00", -- 0x0398
		x"00",x"00",x"01",x"03",x"01",x"00",x"00",x"08", -- 0x03A0
		x"08",x"00",x"00",x"00",x"00",x"60",x"00",x"00", -- 0x03A8
		x"00",x"04",x"92",x"1E",x"8B",x"07",x"0F",x"04", -- 0x03B0
		x"00",x"00",x"00",x"08",x"0C",x"02",x"00",x"00", -- 0x03B8
		x"EE",x"47",x"07",x"01",x"C3",x"70",x"79",x"3B", -- 0x03C0
		x"01",x"80",x"C0",x"C1",x"E3",x"FF",x"FF",x"FF", -- 0x03C8
		x"19",x"3E",x"3F",x"DF",x"57",x"E6",x"E4",x"F0", -- 0x03D0
		x"5C",x"06",x"0E",x"03",x"03",x"85",x"C0",x"F8", -- 0x03D8
		x"3F",x"1F",x"0C",x"83",x"06",x"00",x"80",x"CE", -- 0x03E0
		x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03E8
		x"F7",x"AB",x"13",x"21",x"12",x"05",x"0F",x"06", -- 0x03F0
		x"02",x"0D",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03F8
		x"EE",x"47",x"07",x"01",x"C3",x"70",x"39",x"1F", -- 0x0400
		x"03",x"00",x"81",x"C3",x"F7",x"FF",x"FF",x"FF", -- 0x0408
		x"19",x"3E",x"3F",x"DF",x"57",x"EA",x"C0",x"80", -- 0x0410
		x"84",x"C6",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0418
		x"9F",x"C3",x"6D",x"9F",x"97",x"8E",x"40",x"29", -- 0x0420
		x"1F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0428
		x"CE",x"B3",x"37",x"87",x"2F",x"FF",x"FF",x"FF", -- 0x0430
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0438
		x"DB",x"BC",x"37",x"74",x"B8",x"56",x"E9",x"D4", -- 0x0440
		x"CC",x"A7",x"43",x"82",x"41",x"A5",x"9A",x"EC", -- 0x0448
		x"5D",x"66",x"2B",x"37",x"5B",x"39",x"D5",x"AB", -- 0x0450
		x"DD",x"45",x"77",x"D3",x"62",x"55",x"DB",x"E7", -- 0x0458
		x"85",x"D3",x"6D",x"8E",x"34",x"17",x"D9",x"A4", -- 0x0460
		x"56",x"AA",x"40",x"14",x"66",x"99",x"85",x"4E", -- 0x0468
		x"C9",x"23",x"25",x"C9",x"8A",x"47",x"65",x"42", -- 0x0470
		x"2A",x"51",x"C4",x"4A",x"6D",x"37",x"19",x"BB", -- 0x0478
		x"3F",x"9F",x"6C",x"D3",x"EA",x"AD",x"B2",x"97", -- 0x0480
		x"DF",x"85",x"E1",x"4C",x"D0",x"C2",x"75",x"BE", -- 0x0488
		x"F7",x"A3",x"D3",x"61",x"52",x"05",x"89",x"5D", -- 0x0490
		x"6A",x"59",x"1D",x"2D",x"1B",x"06",x"09",x"CF", -- 0x0498
		x"EE",x"47",x"07",x"01",x"C3",x"50",x"69",x"BF", -- 0x04A0
		x"93",x"F8",x"69",x"16",x"62",x"2A",x"BD",x"EF", -- 0x04A8
		x"19",x"3A",x"3D",x"DD",x"57",x"A6",x"C4",x"D0", -- 0x04B0
		x"7C",x"D6",x"26",x"D3",x"E3",x"79",x"34",x"FE", -- 0x04B8
		x"FF",x"FD",x"DF",x"BF",x"FF",x"FD",x"FF",x"FF", -- 0x04C0
		x"FF",x"FF",x"FF",x"DF",x"FF",x"FF",x"FE",x"FF", -- 0x04C8
		x"FF",x"FF",x"EF",x"FD",x"FF",x"7F",x"FB",x"FF", -- 0x04D0
		x"FF",x"FF",x"FF",x"FF",x"3D",x"BF",x"FF",x"FF", -- 0x04D8
		x"FF",x"F7",x"B7",x"FF",x"F6",x"DF",x"FF",x"FF", -- 0x04E0
		x"FF",x"F7",x"FD",x"E7",x"FF",x"FF",x"FF",x"FF", -- 0x04E8
		x"FF",x"FF",x"F3",x"F3",x"F7",x"FF",x"DF",x"AF", -- 0x04F0
		x"FF",x"FB",x"FD",x"E9",x"EF",x"CF",x"E7",x"FF", -- 0x04F8
		x"00",x"02",x"00",x"00",x"21",x"00",x"08",x"01", -- 0x0500
		x"00",x"03",x"01",x"00",x"00",x"02",x"00",x"00", -- 0x0508
		x"FF",x"47",x"0F",x"1F",x"9F",x"BF",x"43",x"A1", -- 0x0510
		x"14",x"80",x"60",x"24",x"06",x"00",x"00",x"00", -- 0x0518
		x"7F",x"3F",x"1F",x"3F",x"21",x"23",x"76",x"64", -- 0x0520
		x"24",x"10",x"00",x"00",x"00",x"18",x"0C",x"00", -- 0x0528
		x"FF",x"FF",x"FF",x"EF",x"9F",x"8F",x"DF",x"13", -- 0x0530
		x"18",x"38",x"38",x"30",x"12",x"42",x"60",x"00", -- 0x0538
		x"7F",x"7F",x"13",x"07",x"07",x"1E",x"10",x"31", -- 0x0540
		x"02",x"63",x"13",x"20",x"04",x"0E",x"00",x"00", -- 0x0548
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"AF", -- 0x0550
		x"9F",x"3F",x"1F",x"9F",x"93",x"C7",x"01",x"10", -- 0x0558
		x"FF",x"FF",x"FF",x"FF",x"FB",x"FD",x"FB",x"F3", -- 0x0560
		x"47",x"21",x"61",x"70",x"00",x"04",x"08",x"00", -- 0x0568
		x"FF",x"FF",x"BF",x"DF",x"C7",x"C7",x"EF",x"FF", -- 0x0570
		x"FF",x"FF",x"FF",x"3F",x"1F",x"1F",x"23",x"00", -- 0x0578
		x"7F",x"3F",x"1F",x"1F",x"1F",x"47",x"4F",x"0F", -- 0x0580
		x"2F",x"07",x"86",x"64",x"39",x"21",x"44",x"02", -- 0x0588
		x"FF",x"DF",x"8F",x"C7",x"DF",x"FF",x"FF",x"FF", -- 0x0590
		x"FF",x"BF",x"CF",x"DF",x"FF",x"FF",x"FF",x"FF", -- 0x0598
		x"FF",x"FF",x"F9",x"FC",x"F4",x"F8",x"FB",x"7F", -- 0x05A0
		x"3F",x"1D",x"39",x"63",x"43",x"A7",x"62",x"00", -- 0x05A8
		x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"FF",x"CF", -- 0x05B0
		x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05B8
		x"00",x"03",x"26",x"08",x"02",x"06",x"0C",x"00", -- 0x05C0
		x"02",x"03",x"01",x"22",x"04",x"12",x"00",x"00", -- 0x05C8
		x"FF",x"FF",x"7F",x"FF",x"5F",x"3F",x"5F",x"2F", -- 0x05D0
		x"7F",x"DB",x"8D",x"89",x"43",x"03",x"03",x"00", -- 0x05D8
		x"00",x"40",x"00",x"01",x"01",x"20",x"00",x"00", -- 0x05E0
		x"04",x"00",x"00",x"40",x"01",x"00",x"02",x"00", -- 0x05E8
		x"00",x"88",x"00",x"00",x"00",x"00",x"08",x"04", -- 0x05F0
		x"00",x"00",x"04",x"00",x"00",x"01",x"08",x"00", -- 0x05F8
		x"00",x"01",x"00",x"40",x"80",x"00",x"04",x"20", -- 0x0600
		x"00",x"00",x"20",x"24",x"06",x"00",x"00",x"00", -- 0x0608
		x"00",x"18",x"00",x"82",x"C0",x"00",x"04",x"04", -- 0x0610
		x"0A",x"00",x"40",x"80",x"00",x"10",x"00",x"02", -- 0x0618
		x"00",x"08",x"00",x"01",x"01",x"00",x"30",x"00", -- 0x0620
		x"01",x"00",x"00",x"20",x"00",x"80",x"00",x"00", -- 0x0628
		x"10",x"18",x"00",x"00",x"80",x"00",x"04",x"00", -- 0x0630
		x"00",x"00",x"08",x"0C",x"00",x"00",x"41",x"00", -- 0x0638
		x"00",x"00",x"20",x"00",x"00",x"44",x"00",x"00", -- 0x0640
		x"00",x"01",x"22",x"A0",x"00",x"00",x"00",x"00", -- 0x0648
		x"00",x"08",x"00",x"00",x"40",x"20",x"00",x"00", -- 0x0650
		x"00",x"21",x"80",x"00",x"00",x"08",x"40",x"00", -- 0x0658
		x"00",x"08",x"00",x"00",x"00",x"00",x"20",x"00", -- 0x0660
		x"06",x"9B",x"27",x"07",x"13",x"00",x"04",x"00", -- 0x0668
		x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"00", -- 0x0670
		x"00",x"04",x"00",x"C0",x"00",x"00",x"00",x"00", -- 0x0678
		x"00",x"10",x"00",x"20",x"00",x"00",x"40",x"00", -- 0x0680
		x"00",x"00",x"00",x"00",x"40",x"00",x"00",x"00", -- 0x0688
		x"00",x"00",x"10",x"00",x"00",x"00",x"00",x"00", -- 0x0690
		x"40",x"06",x"0F",x"07",x"0F",x"05",x"00",x"00", -- 0x0698
		x"FF",x"FF",x"FF",x"FB",x"57",x"01",x"92",x"09", -- 0x06A0
		x"0D",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06B8
		x"FF",x"FF",x"FF",x"FD",x"F8",x"F8",x"F8",x"FC", -- 0x06C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06C8
		x"FF",x"FF",x"DF",x"0F",x"1F",x"D7",x"6F",x"FD", -- 0x06D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06D8
		x"FD",x"BF",x"FF",x"FD",x"FF",x"E7",x"F4",x"FF", -- 0x06E0
		x"CF",x"DF",x"FB",x"F9",x"BD",x"FF",x"FF",x"FF", -- 0x06E8
		x"FF",x"4F",x"CF",x"DF",x"FE",x"7F",x"7F",x"FB", -- 0x06F0
		x"FF",x"FF",x"EF",x"F7",x"ED",x"FB",x"E7",x"FF", -- 0x06F8
		x"FF",x"FB",x"FC",x"F9",x"FF",x"FF",x"DB",x"C7", -- 0x0700
		x"4C",x"0C",x"08",x"00",x"04",x"36",x"4E",x"04", -- 0x0708
		x"FF",x"FF",x"F7",x"FF",x"FF",x"F7",x"E7",x"31", -- 0x0710
		x"90",x"BE",x"6C",x"42",x"52",x"70",x"00",x"00", -- 0x0718
		x"FF",x"FC",x"FD",x"DF",x"EF",x"EE",x"FE",x"FC", -- 0x0720
		x"FE",x"FE",x"EE",x"F3",x"E3",x"F1",x"F5",x"EF", -- 0x0728
		x"08",x"0C",x"04",x"70",x"D0",x"C6",x"C6",x"4F", -- 0x0730
		x"7B",x"00",x"00",x"80",x"C6",x"CC",x"8C",x"00", -- 0x0738
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0740
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0748
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0750
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0758
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0760
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0768
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0788
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0790
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0800
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0808
		x"08",x"84",x"C0",x"C0",x"C0",x"C0",x"E0",x"E2", -- 0x0810
		x"F0",x"F0",x"F8",x"F8",x"FC",x"FC",x"FE",x"FF", -- 0x0818
		x"80",x"C8",x"C0",x"F0",x"E0",x"F0",x"F8",x"FC", -- 0x0820
		x"FC",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0828
		x"00",x"08",x"04",x"08",x"00",x"20",x"00",x"00", -- 0x0830
		x"00",x"10",x"00",x"02",x"52",x"00",x"00",x"80", -- 0x0838
		x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0840
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0848
		x"80",x"02",x"04",x"00",x"08",x"80",x"00",x"C0", -- 0x0850
		x"C0",x"80",x"06",x"82",x"C4",x"80",x"00",x"80", -- 0x0858
		x"00",x"12",x"10",x"00",x"00",x"00",x"20",x"C0", -- 0x0860
		x"E2",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0868
		x"00",x"00",x"08",x"00",x"00",x"40",x"80",x"40", -- 0x0870
		x"08",x"04",x"10",x"80",x"C0",x"F8",x"FE",x"FF", -- 0x0878
		x"00",x"00",x"13",x"00",x"00",x"00",x"A1",x"80", -- 0x0880
		x"E4",x"F8",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF", -- 0x0888
		x"00",x"88",x"88",x"00",x"00",x"00",x"00",x"02", -- 0x0890
		x"02",x"80",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x0898
		x"00",x"20",x"20",x"01",x"08",x"40",x"61",x"F7", -- 0x08A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08A8
		x"00",x"04",x"20",x"20",x"90",x"80",x"80",x"83", -- 0x08B0
		x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08B8
		x"80",x"E4",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08C8
		x"00",x"82",x"00",x"00",x"80",x"F0",x"FC",x"FE", -- 0x08D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08E8
		x"80",x"D0",x"D4",x"F0",x"E0",x"F5",x"FE",x"FE", -- 0x08F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08F8
		x"89",x"D0",x"F4",x"F8",x"FC",x"FE",x"FF",x"FE", -- 0x0900
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0908
		x"00",x"90",x"10",x"44",x"06",x"80",x"02",x"20", -- 0x0910
		x"20",x"F0",x"F0",x"F4",x"F4",x"FC",x"FE",x"FF", -- 0x0918
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0920
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0928
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0930
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0938
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0940
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0948
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0950
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0958
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0960
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0968
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0978
		x"80",x"88",x"C0",x"F0",x"E0",x"C0",x"E0",x"F4", -- 0x0980
		x"E0",x"F0",x"F2",x"F8",x"F4",x"F8",x"F0",x"F8", -- 0x0988
		x"00",x"08",x"04",x"88",x"80",x"40",x"00",x"00", -- 0x0990
		x"00",x"10",x"00",x"02",x"52",x"00",x"00",x"80", -- 0x0998
		x"F0",x"F8",x"F0",x"FE",x"FC",x"FE",x"FE",x"FD", -- 0x09A0
		x"FE",x"FC",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09A8
		x"80",x"02",x"04",x"00",x"08",x"80",x"00",x"00", -- 0x09B0
		x"00",x"80",x"06",x"82",x"C4",x"80",x"00",x"80", -- 0x09B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09C8
		x"08",x"84",x"C0",x"C0",x"C0",x"C0",x"E0",x"E6", -- 0x09D0
		x"D2",x"E0",x"E0",x"F8",x"F4",x"F0",x"F8",x"F9", -- 0x09D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09E8
		x"F8",x"F4",x"FC",x"F8",x"FC",x"F8",x"FA",x"FE", -- 0x09F0
		x"FC",x"FE",x"FC",x"FE",x"FF",x"FE",x"FE",x"FF", -- 0x09F8
		x"F9",x"F0",x"FC",x"FC",x"FE",x"FE",x"FF",x"FF", -- 0x0A00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A08
		x"00",x"90",x"10",x"44",x"06",x"80",x"02",x"20", -- 0x0A10
		x"20",x"F0",x"F0",x"F4",x"F4",x"FC",x"FE",x"FF", -- 0x0A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A28
		x"F0",x"FA",x"F4",x"F0",x"E8",x"F0",x"E0",x"F0", -- 0x0A30
		x"F8",x"F8",x"F6",x"F2",x"E0",x"E0",x"F0",x"F0", -- 0x0A38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A58
		x"C2",x"C6",x"C4",x"C4",x"C4",x"C4",x"CC",x"C9", -- 0x0A60
		x"C9",x"D9",x"D1",x"D1",x"D3",x"D3",x"D3",x"F3", -- 0x0A68
		x"70",x"60",x"60",x"E7",x"E7",x"C7",x"C7",x"C7", -- 0x0A70
		x"C1",x"CD",x"CD",x"8D",x"81",x"81",x"81",x"81", -- 0x0A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x0A80
		x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A88
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF", -- 0x0A90
		x"FF",x"FF",x"07",x"F7",x"F7",x"F0",x"FE",x"FE", -- 0x0A98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"FF", -- 0x0AA8
		x"FE",x"FF",x"F7",x"F7",x"F7",x"F7",x"F7",x"F7", -- 0x0AB0
		x"F7",x"F7",x"F7",x"F7",x"F7",x"F7",x"F0",x"FE", -- 0x0AB8
		x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"E6",x"F7", -- 0x0AC0
		x"F7",x"F7",x"F7",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x0AC8
		x"FE",x"FF",x"F7",x"FF",x"FF",x"FF",x"07",x"F7", -- 0x0AD0
		x"F7",x"F7",x"F7",x"F7",x"F7",x"F7",x"F0",x"FE", -- 0x0AD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"6F", -- 0x0AE0
		x"4F",x"43",x"47",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x0AE8
		x"FE",x"FF",x"DF",x"DF",x"DF",x"FF",x"FF",x"FF", -- 0x0AF0
		x"FF",x"FF",x"FF",x"1F",x"DF",x"C0",x"FE",x"FE", -- 0x0AF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"EF", -- 0x0B00
		x"EF",x"EF",x"FF",x"BF",x"BF",x"80",x"FF",x"FF", -- 0x0B08
		x"FE",x"FF",x"FD",x"FD",x"FD",x"FD",x"FF",x"EF", -- 0x0B10
		x"EF",x"EF",x"FF",x"FF",x"FF",x"00",x"FE",x"FE", -- 0x0B18
		x"FF",x"FF",x"BC",x"B8",x"B8",x"B8",x"88",x"F8", -- 0x0B20
		x"FF",x"C1",x"81",x"81",x"81",x"83",x"FF",x"FF", -- 0x0B28
		x"FF",x"FF",x"5F",x"5F",x"5F",x"5F",x"5F",x"DF", -- 0x0B30
		x"DF",x"DF",x"DF",x"DF",x"DF",x"C3",x"FF",x"FF", -- 0x0B38
		x"FF",x"CC",x"88",x"88",x"98",x"F8",x"FF",x"BF", -- 0x0B40
		x"BF",x"BF",x"81",x"FF",x"DF",x"DF",x"DF",x"C0", -- 0x0B48
		x"FF",x"7F",x"5F",x"5F",x"5F",x"C3",x"FF",x"87", -- 0x0B50
		x"07",x"07",x"0F",x"F1",x"E1",x"E1",x"E3",x"3F", -- 0x0B58
		x"FF",x"FF",x"DF",x"DF",x"DF",x"DF",x"DF",x"DF", -- 0x0B60
		x"DF",x"C3",x"FF",x"FF",x"EF",x"EF",x"EF",x"E0", -- 0x0B68
		x"FF",x"8F",x"0F",x"0F",x"09",x"01",x"01",x"01", -- 0x0B70
		x"11",x"F3",x"FF",x"DF",x"DF",x"DF",x"C7",x"FF", -- 0x0B78
		x"FF",x"FF",x"BF",x"BF",x"87",x"FC",x"F8",x"F0", -- 0x0B80
		x"E0",x"E0",x"E1",x"F3",x"FF",x"BF",x"87",x"FF", -- 0x0B88
		x"FF",x"F3",x"E1",x"C1",x"81",x"83",x"07",x"4F", -- 0x0B90
		x"7F",x"E7",x"C3",x"83",x"03",x"07",x"0F",x"9F", -- 0x0B98
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA8
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC8
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0BD0
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0BD8
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BE8
		x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0BF0
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0BF8
		x"5F",x"BE",x"F7",x"54",x"68",x"1E",x"2F",x"96", -- 0x0C00
		x"8E",x"C7",x"C3",x"E1",x"F8",x"F9",x"F2",x"F1", -- 0x0C08
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"D5",x"EB", -- 0x0C10
		x"FF",x"77",x"77",x"D3",x"62",x"F5",x"FF",x"27", -- 0x0C18
		x"FC",x"FC",x"9E",x"8F",x"9F",x"FF",x"FF",x"FF", -- 0x0C20
		x"FB",x"F1",x"C3",x"27",x"7F",x"FF",x"F7",x"8F", -- 0x0C28
		x"77",x"3B",x"53",x"09",x"82",x"C1",x"E7",x"E5", -- 0x0C30
		x"E2",x"CF",x"D4",x"8A",x"2D",x"3F",x"99",x"9B", -- 0x0C38
		x"CF",x"FF",x"FF",x"FF",x"FF",x"F7",x"F7",x"6F", -- 0x0C40
		x"1F",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C48
		x"97",x"DB",x"B3",x"81",x"C2",x"C1",x"E7",x"E1", -- 0x0C50
		x"C2",x"E1",x"F1",x"F1",x"F8",x"F9",x"F8",x"FC", -- 0x0C58
		x"3F",x"1F",x"8D",x"C0",x"E2",x"FF",x"FF",x"7F", -- 0x0C60
		x"1F",x"3D",x"3D",x"9B",x"DF",x"DF",x"FE",x"BC", -- 0x0C68
		x"F7",x"AB",x"D3",x"E1",x"52",x"45",x"07",x"82", -- 0x0C70
		x"D9",x"FD",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x0C78
		x"90",x"30",x"61",x"63",x"FF",x"F3",x"F0",x"81", -- 0x0C80
		x"87",x"0F",x"9F",x"BE",x"BC",x"60",x"C1",x"87", -- 0x0C88
		x"79",x"F3",x"F3",x"E7",x"C3",x"87",x"4F",x"DF", -- 0x0C90
		x"DF",x"1F",x"3C",x"38",x"38",x"71",x"E1",x"F7", -- 0x0C98
		x"7F",x"FC",x"C9",x"33",x"CE",x"F1",x"FC",x"FF", -- 0x0CA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CA8
		x"BF",x"FF",x"9C",x"01",x"61",x"73",x"BF",x"CF", -- 0x0CB0
		x"E0",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0CC0
		x"00",x"00",x"00",x"00",x"0F",x"3F",x"FF",x"FF", -- 0x0CC8
		x"17",x"0B",x"13",x"01",x"02",x"01",x"07",x"01", -- 0x0CD0
		x"02",x"01",x"01",x"01",x"80",x"E0",x"F8",x"FC", -- 0x0CD8
		x"1F",x"8F",x"CF",x"CE",x"C7",x"E7",x"E7",x"F3", -- 0x0CE0
		x"33",x"39",x"19",x"99",x"EC",x"EC",x"3C",x"1E", -- 0x0CE8
		x"FE",x"FF",x"77",x"73",x"73",x"E3",x"E3",x"F6", -- 0x0CF0
		x"F7",x"F3",x"BB",x"9D",x"DC",x"DC",x"CE",x"6E", -- 0x0CF8
		x"8E",x"86",x"C3",x"C3",x"E6",x"E6",x"F6",x"F3", -- 0x0D00
		x"F9",x"78",x"7C",x"1C",x"0E",x"8E",x"C7",x"E3", -- 0x0D08
		x"7C",x"3D",x"7B",x"BA",x"72",x"74",x"38",x"18", -- 0x0D10
		x"19",x"99",x"9C",x"CC",x"4D",x"47",x"26",x"26", -- 0x0D18
		x"F3",x"F9",x"F8",x"FD",x"FF",x"FE",x"FE",x"FF", -- 0x0D20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D28
		x"E9",x"F2",x"CD",x"03",x"03",x"01",x"01",x"03", -- 0x0D30
		x"03",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D38
		x"FF",x"FC",x"FD",x"DF",x"EF",x"EE",x"FE",x"FC", -- 0x0D40
		x"FE",x"FE",x"EE",x"F7",x"E2",x"F7",x"FF",x"FF", -- 0x0D48
		x"08",x"04",x"04",x"70",x"50",x"86",x"C3",x"49", -- 0x0D50
		x"3B",x"20",x"08",x"80",x"38",x"FF",x"FF",x"FF", -- 0x0D58
		x"77",x"7F",x"BB",x"BD",x"DF",x"CE",x"E7",x"E7", -- 0x0D60
		x"FF",x"FF",x"FF",x"79",x"7C",x"7C",x"3E",x"3F", -- 0x0D68
		x"FF",x"FF",x"FF",x"F3",x"F3",x"F9",x"7D",x"38", -- 0x0D70
		x"BC",x"BE",x"DF",x"CF",x"FF",x"FF",x"7F",x"7F", -- 0x0D78
		x"9E",x"F7",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D80
		x"FF",x"1F",x"CF",x"FF",x"FF",x"FE",x"FC",x"F8", -- 0x0D88
		x"6F",x"E7",x"E7",x"EF",x"F7",x"F3",x"FB",x"F9", -- 0x0D90
		x"FC",x"FF",x"DF",x"8F",x"CF",x"F7",x"FB",x"FB", -- 0x0D98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DD0
		x"FF",x"FF",x"FF",x"DF",x"EF",x"E7",x"F7",x"F3", -- 0x0DD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E60
		x"91",x"A0",x"50",x"20",x"10",x"08",x"00",x"00", -- 0x0E68
		x"00",x"00",x"80",x"40",x"64",x"28",x"54",x"08", -- 0x0E70
		x"04",x"80",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E78
		x"00",x"00",x"08",x"04",x"06",x"02",x"05",x"00", -- 0x0E80
		x"10",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E88
		x"00",x"00",x"00",x"00",x"40",x"80",x"42",x"81", -- 0x0E90
		x"41",x"20",x"01",x"00",x"04",x"02",x"00",x"00", -- 0x0E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0ED8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF8
		x"80",x"C0",x"E0",x"E0",x"E0",x"E6",x"EE",x"7C", -- 0x1000
		x"70",x"B8",x"B8",x"BA",x"DE",x"5C",x"AC",x"F6", -- 0x1008
		x"00",x"00",x"00",x"08",x"00",x"00",x"00",x"00", -- 0x1010
		x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1018
		x"36",x"1B",x"1D",x"3F",x"7F",x"6F",x"CD",x"C7", -- 0x1020
		x"85",x"CF",x"DF",x"FB",x"F1",x"61",x"61",x"38", -- 0x1028
		x"00",x"80",x"80",x"C0",x"D0",x"F0",x"E0",x"C0", -- 0x1030
		x"80",x"98",x"F0",x"E0",x"E4",x"E8",x"F0",x"E6", -- 0x1038
		x"7F",x"BB",x"B8",x"99",x"BE",x"FD",x"DA",x"CC", -- 0x1040
		x"5C",x"EC",x"FF",x"F7",x"76",x"3F",x"FF",x"FF", -- 0x1048
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"76",x"3C", -- 0x1050
		x"78",x"F8",x"F8",x"38",x"3B",x"FE",x"FC",x"FC", -- 0x1058
		x"00",x"80",x"C0",x"D0",x"F0",x"E0",x"F0",x"7C", -- 0x1060
		x"78",x"38",x"38",x"3A",x"1C",x"1F",x"CE",x"C6", -- 0x1068
		x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00", -- 0x1070
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1078
		x"EF",x"FF",x"F7",x"E3",x"F7",x"FF",x"F3",x"79", -- 0x1080
		x"7B",x"7F",x"7D",x"38",x"3C",x"BD",x"9D",x"FF", -- 0x1088
		x"40",x"E0",x"80",x"C0",x"C0",x"C0",x"E8",x"F8", -- 0x1090
		x"E0",x"C0",x"E0",x"E0",x"C0",x"C4",x"C8",x"D8", -- 0x1098
		x"66",x"26",x"16",x"1B",x"1B",x"3D",x"26",x"C7", -- 0x10A0
		x"E3",x"E3",x"E3",x"E7",x"E5",x"FD",x"F8",x"F0", -- 0x10A8
		x"70",x"FC",x"F0",x"E0",x"70",x"E0",x"44",x"4C", -- 0x10B0
		x"78",x"30",x"F0",x"B0",x"B0",x"B2",x"9A",x"8C", -- 0x10B8
		x"F8",x"D8",x"CD",x"FF",x"6E",x"37",x"3F",x"9B", -- 0x10C0
		x"DF",x"FD",x"EF",x"7F",x"3F",x"3F",x"1B",x"18", -- 0x10C8
		x"76",x"F7",x"BB",x"7B",x"7B",x"FD",x"DD",x"9C", -- 0x10D0
		x"9F",x"EF",x"DF",x"FB",x"31",x"99",x"FD",x"FC", -- 0x10D8
		x"CF",x"C7",x"69",x"79",x"78",x"99",x"9B",x"8F", -- 0x10E0
		x"CE",x"E7",x"EF",x"FB",x"F1",x"E3",x"F7",x"FE", -- 0x10E8
		x"F8",x"F1",x"FB",x"FE",x"BE",x"FE",x"DF",x"7F", -- 0x10F0
		x"6F",x"37",x"3B",x"9F",x"9E",x"FF",x"F7",x"E3", -- 0x10F8
		x"3B",x"1E",x"3C",x"7C",x"FE",x"FF",x"FF",x"FB", -- 0x1100
		x"F9",x"71",x"39",x"BF",x"FE",x"BC",x"3F",x"7F", -- 0x1108
		x"F9",x"78",x"3C",x"1D",x"3B",x"DB",x"1B",x"19", -- 0x1110
		x"CC",x"8D",x"FD",x"FD",x"7D",x"E4",x"C4",x"E6", -- 0x1118
		x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00", -- 0x1120
		x"00",x"00",x"1C",x"3F",x"1F",x"0F",x"1F",x"1F", -- 0x1128
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1130
		x"00",x"00",x"00",x"F0",x"F8",x"FC",x"FE",x"FE", -- 0x1138
		x"30",x"60",x"80",x"80",x"C0",x"C0",x"60",x"61", -- 0x1140
		x"37",x"7F",x"FF",x"FF",x"FF",x"FF",x"F8",x"E0", -- 0x1148
		x"7F",x"3F",x"3F",x"3F",x"3F",x"3D",x"39",x"F0", -- 0x1150
		x"F8",x"F8",x"FE",x"FE",x"FF",x"FF",x"1F",x"0F", -- 0x1158
		x"0F",x"9F",x"7F",x"FF",x"FF",x"FF",x"FE",x"F9", -- 0x1160
		x"E3",x"C7",x"8F",x"9F",x"3F",x"7C",x"E0",x"C0", -- 0x1168
		x"C7",x"F1",x"F9",x"FC",x"FE",x"FF",x"0F",x"F7", -- 0x1170
		x"FB",x"F9",x"FD",x"FE",x"8E",x"03",x"00",x"00", -- 0x1178
		x"C0",x"00",x"03",x"07",x"0F",x"0F",x"1F",x"3F", -- 0x1180
		x"7F",x"FF",x"FF",x"F7",x"E7",x"CF",x"9F",x"9F", -- 0x1188
		x"08",x"3C",x"FC",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x1190
		x"F7",x"F3",x"F9",x"FC",x"FE",x"FF",x"FF",x"0F", -- 0x1198
		x"1D",x"33",x"67",x"4F",x"DF",x"BE",x"3C",x"39", -- 0x11A0
		x"73",x"CF",x"9F",x"1C",x"38",x"78",x"F0",x"F0", -- 0x11A8
		x"F9",x"FE",x"FF",x"83",x"38",x"7C",x"FF",x"FF", -- 0x11B0
		x"FF",x"E3",x"00",x"00",x"3C",x"7F",x"FF",x"FF", -- 0x11B8
		x"D9",x"DF",x"8F",x"87",x"8F",x"8F",x"0F",x"0E", -- 0x11C0
		x"1E",x"1C",x"3C",x"38",x"38",x"38",x"70",x"70", -- 0x11C8
		x"FF",x"F8",x"F0",x"E0",x"C0",x"C0",x"E1",x"F3", -- 0x11D0
		x"7F",x"3F",x"3F",x"7F",x"7F",x"FF",x"FF",x"FF", -- 0x11D8
		x"70",x"F0",x"E1",x"E1",x"E3",x"C3",x"C7",x"C7", -- 0x11E0
		x"C7",x"C7",x"C7",x"C7",x"E3",x"EF",x"CF",x"CE", -- 0x11E8
		x"FE",x"FE",x"F3",x"E3",x"E7",x"CF",x"CF",x"8F", -- 0x11F0
		x"8F",x"1F",x"39",x"3C",x"3E",x"3F",x"B1",x"72", -- 0x11F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1200
		x"0C",x"06",x"03",x"03",x"07",x"0F",x"0F",x"1F", -- 0x1208
		x"08",x"10",x"31",x"73",x"3F",x"3E",x"7C",x"7C", -- 0x1210
		x"F4",x"E6",x"E2",x"C1",x"81",x"83",x"C7",x"E7", -- 0x1218
		x"7E",x"FC",x"F8",x"F0",x"F0",x"F0",x"E1",x"E1", -- 0x1220
		x"E0",x"E0",x"F0",x"99",x"9D",x"9F",x"1D",x"1D", -- 0x1228
		x"6F",x"3E",x"3C",x"78",x"70",x"F1",x"F3",x"F7", -- 0x1230
		x"E7",x"E7",x"EF",x"EF",x"EF",x"DF",x"DF",x"9F", -- 0x1238
		x"3B",x"37",x"37",x"77",x"6E",x"6E",x"6E",x"6E", -- 0x1240
		x"EE",x"EE",x"E4",x"F1",x"F9",x"EE",x"ED",x"EC", -- 0x1248
		x"9E",x"9E",x"BC",x"3C",x"78",x"F8",x"F8",x"F0", -- 0x1250
		x"B0",x"60",x"E0",x"C0",x"C1",x"C3",x"E3",x"E7", -- 0x1258
		x"EC",x"CC",x"DC",x"9E",x"9E",x"3E",x"7E",x"7E", -- 0x1260
		x"7F",x"7D",x"FC",x"FC",x"78",x"78",x"78",x"78", -- 0x1268
		x"67",x"37",x"0F",x"06",x"06",x"0C",x"0C",x"0C", -- 0x1270
		x"0C",x"CC",x"78",x"19",x"1B",x"3B",x"F3",x"E7", -- 0x1278
		x"31",x"31",x"18",x"86",x"C3",x"C1",x"E1",x"FB", -- 0x1280
		x"9F",x"8F",x"8F",x"8F",x"8F",x"8F",x"86",x"86", -- 0x1288
		x"E2",x"E4",x"F9",x"D9",x"D9",x"E3",x"D7",x"B7", -- 0x1290
		x"FF",x"9F",x"6E",x"6E",x"9C",x"3C",x"D8",x"D8", -- 0x1298
		x"8F",x"0E",x"1E",x"1B",x"37",x"36",x"36",x"36", -- 0x12A0
		x"7F",x"7B",x"79",x"37",x"36",x"32",x"10",x"1B", -- 0x12A8
		x"38",x"78",x"70",x"30",x"60",x"E0",x"E1",x"E1", -- 0x12B0
		x"E1",x"61",x"31",x"70",x"70",x"7D",x"3F",x"37", -- 0x12B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12D0
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x12D8
		x"00",x"00",x"10",x"08",x"00",x"00",x"00",x"00", -- 0x12E0
		x"00",x"40",x"00",x"00",x"01",x"00",x"00",x"00", -- 0x12E8
		x"00",x"08",x"04",x"06",x"03",x"01",x"00",x"01", -- 0x12F0
		x"03",x"43",x"F7",x"3F",x"1F",x"0F",x"0F",x"0F", -- 0x12F8
		x"00",x"00",x"00",x"00",x"00",x"03",x"00",x"00", -- 0x1300
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1308
		x"0F",x"1E",x"1E",x"1E",x"3E",x"3E",x"FC",x"3C", -- 0x1310
		x"38",x"78",x"78",x"7C",x"7C",x"78",x"38",x"38", -- 0x1318
		x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1320
		x"04",x"03",x"03",x"03",x"03",x"07",x"03",x"03", -- 0x1328
		x"71",x"F3",x"73",x"7B",x"6F",x"E7",x"E7",x"F7", -- 0x1330
		x"C7",x"C6",x"8E",x"8E",x"EE",x"AE",x"9E",x"9E", -- 0x1338
		x"03",x"03",x"03",x"17",x"3F",x"1F",x"0F",x"07", -- 0x1340
		x"07",x"07",x"03",x"03",x"03",x"03",x"33",x"39", -- 0x1348
		x"EF",x"FF",x"BF",x"9F",x"DF",x"FF",x"3F",x"3F", -- 0x1350
		x"3F",x"3F",x"3F",x"1F",x"9F",x"9F",x"8F",x"CF", -- 0x1358
		x"1F",x"0F",x"07",x"23",x"3F",x"0F",x"07",x"07", -- 0x1360
		x"07",x"07",x"03",x"03",x"13",x"1F",x"03",x"03", -- 0x1368
		x"CF",x"CF",x"E7",x"C7",x"C7",x"8E",x"8E",x"8C", -- 0x1370
		x"0C",x"1C",x"1C",x"DE",x"7E",x"1F",x"1F",x"8F", -- 0x1378
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1380
		x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1388
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1390
		x"00",x"80",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x1398
		x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00", -- 0x13A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F8
		x"7B",x"BF",x"3E",x"7F",x"76",x"FE",x"7D",x"5C", -- 0x1400
		x"CE",x"FD",x"FC",x"BC",x"99",x"F8",x"F9",x"39", -- 0x1408
		x"1C",x"3C",x"3E",x"79",x"78",x"38",x"B8",x"FC", -- 0x1410
		x"3E",x"72",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x1418
		x"3F",x"67",x"63",x"F3",x"EB",x"C7",x"F7",x"9D", -- 0x1420
		x"8D",x"1D",x"0F",x"8F",x"FF",x"7D",x"1B",x"36", -- 0x1428
		x"E0",x"F0",x"F8",x"FC",x"FC",x"F8",x"C8",x"C0", -- 0x1430
		x"E0",x"E0",x"F0",x"F0",x"E0",x"80",x"80",x"00", -- 0x1438
		x"F6",x"AC",x"5C",x"DC",x"B8",x"B0",x"BC",x"7C", -- 0x1440
		x"7C",x"F8",x"F8",x"D8",x"80",x"00",x"00",x"00", -- 0x1448
		x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00", -- 0x1450
		x"00",x"00",x"00",x"10",x"08",x"00",x"00",x"00", -- 0x1458
		x"9E",x"BC",x"7E",x"7F",x"DF",x"1D",x"39",x"7F", -- 0x1460
		x"F7",x"E7",x"EF",x"FF",x"FF",x"5E",x"1E",x"38", -- 0x1468
		x"F7",x"76",x"E6",x"E6",x"F7",x"FF",x"CF",x"CF", -- 0x1470
		x"9E",x"9E",x"FF",x"3F",x"1D",x"3C",x"78",x"F9", -- 0x1478
		x"F0",x"F1",x"E3",x"E6",x"EC",x"CC",x"C9",x"99", -- 0x1480
		x"13",x"33",x"27",x"66",x"CE",x"CE",x"9C",x"9C", -- 0x1488
		x"C8",x"91",x"11",x"21",x"63",x"C7",x"CF",x"8F", -- 0x1490
		x"9E",x"1C",x"18",x"18",x"30",x"30",x"30",x"60", -- 0x1498
		x"3C",x"FE",x"BB",x"F1",x"FB",x"FF",x"FF",x"CF", -- 0x14A0
		x"8E",x"9C",x"9C",x"FC",x"F9",x"F9",x"FF",x"CF", -- 0x14A8
		x"F0",x"F1",x"FB",x"9F",x"9F",x"3B",x"3B",x"FF", -- 0x14B0
		x"FF",x"7F",x"FF",x"FE",x"FE",x"FE",x"FD",x"FD", -- 0x14B8
		x"1C",x"BC",x"BD",x"F9",x"F9",x"F1",x"F3",x"E3", -- 0x14C0
		x"E7",x"C6",x"4C",x"6B",x"3F",x"1F",x"BE",x"F6", -- 0x14C8
		x"EE",x"DE",x"DE",x"DC",x"FC",x"FC",x"BC",x"3C", -- 0x14D0
		x"7E",x"7E",x"78",x"F8",x"F8",x"F8",x"F0",x"70", -- 0x14D8
		x"FC",x"9F",x"BF",x"3C",x"3C",x"79",x"79",x"7D", -- 0x14E0
		x"7F",x"F3",x"F3",x"F3",x"F7",x"FF",x"FF",x"CF", -- 0x14E8
		x"F0",x"E0",x"E0",x"E0",x"E0",x"F0",x"F8",x"F8", -- 0x14F0
		x"E0",x"E0",x"C0",x"E0",x"E0",x"C0",x"80",x"00", -- 0x14F8
		x"CE",x"9E",x"1E",x"1E",x"3C",x"3E",x"7C",x"78", -- 0x1500
		x"F8",x"F0",x"F0",x"E0",x"E0",x"C0",x"C0",x"00", -- 0x1508
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1510
		x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00", -- 0x1518
		x"EE",x"EE",x"EE",x"E7",x"F7",x"C7",x"C7",x"C7", -- 0x1520
		x"C7",x"C7",x"C3",x"E3",x"E1",x"E1",x"F0",x"F1", -- 0x1528
		x"31",x"30",x"38",x"38",x"38",x"3C",x"1E",x"9E", -- 0x1530
		x"8F",x"DF",x"EF",x"E7",x"E3",x"F0",x"F8",x"FE", -- 0x1538
		x"70",x"70",x"38",x"38",x"38",x"3C",x"1C",x"1E", -- 0x1540
		x"0E",x"0F",x"8F",x"8F",x"87",x"8F",x"DF",x"D9", -- 0x1548
		x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"1F",x"0F", -- 0x1550
		x"13",x"21",x"C0",x"C0",x"E1",x"F1",x"FF",x"FF", -- 0x1558
		x"F0",x"F0",x"78",x"38",x"1C",x"9F",x"CF",x"73", -- 0x1560
		x"39",x"3C",x"BE",x"5F",x"4F",x"67",x"33",x"1D", -- 0x1568
		x"FF",x"FF",x"7F",x"1D",x"01",x"00",x"C3",x"FF", -- 0x1570
		x"FF",x"FF",x"7C",x"3E",x"87",x"FF",x"FF",x"FF", -- 0x1578
		x"9F",x"9F",x"CF",x"E7",x"F3",x"F0",x"FC",x"7F", -- 0x1580
		x"3F",x"1F",x"3F",x"3F",x"67",x"E3",x"C0",x"C0", -- 0x1588
		x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"0F", -- 0x1590
		x"9F",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"0F", -- 0x1598
		x"40",x"60",x"7C",x"3F",x"9F",x"8F",x"C7",x"E1", -- 0x15A0
		x"F8",x"FE",x"FF",x"FF",x"FF",x"7F",x"FF",x"EF", -- 0x15A8
		x"0F",x"0F",x"1F",x"9F",x"FF",x"FF",x"FF",x"FF", -- 0x15B0
		x"F7",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"CF", -- 0x15B8
		x"C0",x"F0",x"FF",x"FF",x"FF",x"FF",x"7F",x"37", -- 0x15C0
		x"21",x"60",x"40",x"40",x"80",x"80",x"60",x"30", -- 0x15C8
		x"6F",x"DF",x"FF",x"FF",x"FE",x"FE",x"F8",x"F8", -- 0x15D0
		x"F0",x"21",x"31",x"3B",x"3F",x"1F",x"3F",x"7E", -- 0x15D8
		x"1F",x"1F",x"0F",x"07",x"03",x"00",x"00",x"00", -- 0x15E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15E8
		x"FF",x"FF",x"FE",x"FC",x"FC",x"18",x"10",x"00", -- 0x15F0
		x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"00", -- 0x15F8
		x"1B",x"7F",x"B6",x"F6",x"73",x"FF",x"79",x"3D", -- 0x1600
		x"36",x"36",x"36",x"37",x"3B",x"1D",x"1E",x"8F", -- 0x1608
		x"71",x"F1",x"78",x"78",x"7F",x"7F",x"F7",x"E1", -- 0x1610
		x"E1",x"E1",x"E1",x"60",x"F0",x"F0",x"78",x"7B", -- 0x1618
		x"9E",x"F6",x"CE",x"8F",x"8F",x"8F",x"87",x"87", -- 0x1620
		x"C7",x"DD",x"F9",x"F1",x"E0",x"D6",x"BF",x"B9", -- 0x1628
		x"DE",x"DC",x"5C",x"5C",x"6E",x"6E",x"27",x"B7", -- 0x1630
		x"B7",x"97",x"D7",x"DB",x"DF",x"CD",x"EC",x"FE", -- 0x1638
		x"1F",x"3F",x"3E",x"38",x"7C",x"7C",x"3C",x"3E", -- 0x1640
		x"3E",x"3E",x"1F",x"9F",x"8F",x"CF",x"C6",x"E4", -- 0x1648
		x"63",x"71",x"3F",x"3F",x"1C",x"18",x"0D",x"0F", -- 0x1650
		x"0F",x"46",x"E0",x"C2",x"83",x"03",x"0B",x"5B", -- 0x1658
		x"EC",x"ED",x"EF",x"F7",x"FF",x"F8",x"FC",x"EF", -- 0x1660
		x"6F",x"6F",x"6E",x"66",x"77",x"37",x"37",x"3B", -- 0x1668
		x"E7",x"EF",x"DF",x"FB",x"F0",x"E0",x"E0",x"F0", -- 0x1670
		x"F0",x"F8",x"F8",x"78",x"3C",x"9C",x"9E",x"BE", -- 0x1678
		x"CF",x"0F",x"8D",x"84",x"80",x"C3",x"E7",x"FE", -- 0x1680
		x"FE",x"FC",x"F0",x"F0",x"F0",x"78",x"7C",x"3E", -- 0x1688
		x"EF",x"EE",x"EE",x"EF",x"E7",x"77",x"77",x"E3", -- 0x1690
		x"F3",x"FD",x"7C",x"38",x"38",x"1C",x"0E",x"43", -- 0x1698
		x"7F",x"FF",x"FF",x"7F",x"27",x"01",x"00",x"00", -- 0x16A0
		x"01",x"03",x"03",x"00",x"00",x"00",x"00",x"00", -- 0x16A8
		x"E7",x"C7",x"87",x"83",x"C1",x"E3",x"E7",x"F7", -- 0x16B0
		x"FB",x"FF",x"7F",x"0F",x"03",x"0D",x"0E",x"06", -- 0x16B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16C0
		x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00", -- 0x16C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D8
		x"01",x"03",x"03",x"03",x"1B",x"1F",x"3F",x"07", -- 0x16E0
		x"07",x"07",x"07",x"07",x"07",x"03",x"01",x"03", -- 0x16E8
		x"3F",x"3F",x"FF",x"FF",x"1E",x"1F",x"1F",x"BF", -- 0x16F0
		x"FC",x"8E",x"8E",x"DF",x"E7",x"E7",x"CF",x"FF", -- 0x16F8
		x"03",x"03",x"03",x"1B",x"3F",x"3F",x"17",x"07", -- 0x1700
		x"07",x"07",x"07",x"07",x"07",x"03",x"03",x"01", -- 0x1708
		x"FF",x"FF",x"9F",x"FF",x"FF",x"3F",x"3F",x"3F", -- 0x1710
		x"3F",x"3F",x"3F",x"9F",x"9F",x"9F",x"8F",x"CF", -- 0x1718
		x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"00", -- 0x1720
		x"00",x"00",x"01",x"03",x"06",x"00",x"00",x"00", -- 0x1728
		x"FE",x"DE",x"9E",x"FE",x"EE",x"CE",x"E6",x"EF", -- 0x1730
		x"FF",x"F7",x"E7",x"63",x"77",x"7F",x"7F",x"7F", -- 0x1738
		x"00",x"06",x"07",x"03",x"01",x"00",x"00",x"00", -- 0x1740
		x"00",x"00",x"01",x"03",x"00",x"00",x"00",x"01", -- 0x1748
		x"18",x"38",x"78",x"FF",x"FF",x"7E",x"78",x"78", -- 0x1750
		x"3C",x"7C",x"FE",x"3E",x"1E",x"1E",x"7E",x"DF", -- 0x1758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1760
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1768
		x"CF",x"0F",x"0F",x"07",x"07",x"07",x"07",x"03", -- 0x1770
		x"03",x"01",x"03",x"02",x"06",x"04",x"08",x"00", -- 0x1778
		x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00", -- 0x1780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1798
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17C0
		x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00", -- 0x17C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D8
		x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00", -- 0x17E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17F0
		x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x17F8
		x"00",x"00",x"00",x"08",x"08",x"00",x"00",x"00", -- 0x1800
		x"00",x"00",x"00",x"20",x"00",x"00",x"01",x"00", -- 0x1808
		x"00",x"01",x"00",x"40",x"00",x"02",x"0C",x"04", -- 0x1810
		x"00",x"10",x"22",x"02",x"01",x"00",x"01",x"00", -- 0x1818
		x"81",x"00",x"00",x"02",x"01",x"84",x"02",x"00", -- 0x1820
		x"02",x"01",x"04",x"01",x"00",x"00",x"41",x"00", -- 0x1828
		x"00",x"81",x"80",x"40",x"00",x"02",x"0C",x"04", -- 0x1830
		x"00",x"00",x"01",x"02",x"05",x"02",x"01",x"00", -- 0x1838
		x"89",x"2C",x"04",x"00",x"00",x"00",x"00",x"00", -- 0x1840
		x"00",x"00",x"00",x"01",x"01",x"00",x"40",x"00", -- 0x1848
		x"00",x"81",x"80",x"40",x"00",x"42",x"2C",x"04", -- 0x1850
		x"10",x"00",x"40",x"40",x"50",x"1A",x"CD",x"00", -- 0x1858
		x"81",x"00",x"00",x"02",x"00",x"07",x"02",x"00", -- 0x1860
		x"02",x"00",x"06",x"00",x"00",x"00",x"00",x"01", -- 0x1868
		x"00",x"81",x"80",x"41",x"01",x"42",x"0C",x"05", -- 0x1870
		x"03",x"40",x"82",x"02",x"05",x"02",x"09",x"00", -- 0x1878
		x"81",x"12",x"40",x"02",x"01",x"10",x"00",x"00", -- 0x1880
		x"00",x"00",x"40",x"00",x"00",x"00",x"09",x"00", -- 0x1888
		x"00",x"81",x"80",x"40",x"00",x"42",x"2C",x"04", -- 0x1890
		x"08",x"10",x"00",x"00",x"02",x"00",x"10",x"00", -- 0x1898
		x"81",x"00",x"02",x"08",x"88",x"80",x"00",x"00", -- 0x18A0
		x"00",x"20",x"50",x"00",x"12",x"00",x"00",x"00", -- 0x18A8
		x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"02", -- 0x18B0
		x"00",x"40",x"00",x"00",x"10",x"04",x"04",x"20", -- 0x18B8
		x"6C",x"D2",x"91",x"10",x"00",x"02",x"08",x"48", -- 0x18C0
		x"44",x"22",x"00",x"10",x"80",x"00",x"00",x"00", -- 0x18C8
		x"50",x"A8",x"45",x"C1",x"03",x"04",x"00",x"00", -- 0x18D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
		x"81",x"00",x"00",x"02",x"80",x"84",x"02",x"00", -- 0x18E0
		x"02",x"21",x"54",x"21",x"00",x"20",x"60",x"11", -- 0x18E8
		x"00",x"84",x"82",x"42",x"00",x"44",x"28",x"04", -- 0x18F0
		x"10",x"00",x"02",x"00",x"00",x"00",x"04",x"00", -- 0x18F8
		x"81",x"00",x"00",x"00",x"80",x"84",x"02",x"04", -- 0x1900
		x"00",x"20",x"50",x"02",x"10",x"00",x"00",x"00", -- 0x1908
		x"00",x"80",x"80",x"40",x"00",x"40",x"20",x"02", -- 0x1910
		x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"00", -- 0x1918
		x"81",x"00",x"40",x"00",x"88",x"94",x"02",x"20", -- 0x1920
		x"00",x"00",x"40",x"00",x"00",x"00",x"10",x"00", -- 0x1928
		x"00",x"80",x"80",x"40",x"00",x"40",x"20",x"00", -- 0x1930
		x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1938
		x"00",x"00",x"08",x"00",x"00",x"00",x"00",x"00", -- 0x1940
		x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1948
		x"00",x"02",x"01",x"02",x"00",x"03",x"06",x"02", -- 0x1950
		x"00",x"00",x"01",x"11",x"01",x"00",x"80",x"10", -- 0x1958
		x"00",x"00",x"00",x"00",x"00",x"02",x"08",x"08", -- 0x1960
		x"44",x"22",x"00",x"11",x"82",x"0C",x"4A",x"64", -- 0x1968
		x"01",x"00",x"01",x"0B",x"03",x"04",x"00",x"00", -- 0x1970
		x"00",x"20",x"24",x"06",x"29",x"4C",x"36",x"0C", -- 0x1978
		x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00", -- 0x1980
		x"00",x"0A",x"00",x"11",x"22",x"34",x"2A",x"04", -- 0x1988
		x"50",x"88",x"05",x"81",x"03",x"04",x"00",x"00", -- 0x1990
		x"00",x"20",x"24",x"06",x"29",x"4C",x"36",x"0C", -- 0x1998
		x"00",x"20",x"00",x"01",x"00",x"00",x"00",x"00", -- 0x19A0
		x"00",x"00",x"00",x"01",x"02",x"04",x"4A",x"64", -- 0x19A8
		x"00",x"00",x"01",x"0B",x"03",x"04",x"00",x"00", -- 0x19B0
		x"00",x"20",x"24",x"06",x"29",x"4C",x"36",x"0C", -- 0x19B8
		x"00",x"00",x"40",x"00",x"00",x"04",x"00",x"00", -- 0x19C0
		x"00",x"00",x"00",x"01",x"02",x"0C",x"4A",x"64", -- 0x19C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"00", -- 0x19D0
		x"00",x"42",x"02",x"02",x"01",x"00",x"80",x"10", -- 0x19D8
		x"80",x"40",x"80",x"00",x"80",x"00",x"58",x"08", -- 0x19E0
		x"04",x"23",x"00",x"10",x"80",x"0C",x"4A",x"64", -- 0x19E8
		x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x19F0
		x"00",x"00",x"08",x"08",x"00",x"00",x"00",x"00", -- 0x19F8
		x"80",x"40",x"88",x"18",x"81",x"02",x"58",x"49", -- 0x1A00
		x"44",x"22",x"00",x"11",x"82",x"0C",x"4A",x"64", -- 0x1A08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A10
		x"02",x"01",x"03",x"02",x"01",x"00",x"80",x"10", -- 0x1A18
		x"01",x"02",x"8F",x"10",x"80",x"02",x"58",x"48", -- 0x1A20
		x"44",x"22",x"00",x"11",x"82",x"0C",x"4A",x"64", -- 0x1A28
		x"00",x"80",x"00",x"40",x"00",x"00",x"08",x"04", -- 0x1A30
		x"00",x"20",x"00",x"00",x"02",x"06",x"82",x"11", -- 0x1A38
		x"80",x"40",x"80",x"00",x"80",x"00",x"59",x"08", -- 0x1A40
		x"04",x"22",x"00",x"11",x"80",x"0C",x"4A",x"64", -- 0x1A48
		x"00",x"00",x"04",x"00",x"00",x"00",x"40",x"00", -- 0x1A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"10", -- 0x1A58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A60
		x"44",x"02",x"00",x"01",x"82",x"00",x"42",x"64", -- 0x1A68
		x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A70
		x"00",x"80",x"00",x"04",x"10",x"24",x"82",x"11", -- 0x1A78
		x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A80
		x"02",x"21",x"D4",x"21",x"00",x"20",x"60",x"10", -- 0x1A88
		x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"00", -- 0x1A90
		x"12",x"09",x"43",x"41",x"00",x"0A",x"CD",x"00", -- 0x1A98
		x"81",x"00",x"00",x"02",x"82",x"85",x"00",x"60", -- 0x1AA0
		x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00", -- 0x1AA8
		x"00",x"01",x"00",x"40",x"00",x"42",x"AC",x"10", -- 0x1AB0
		x"10",x"0A",x"10",x"00",x"00",x"08",x"00",x"00", -- 0x1AB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"00", -- 0x1AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC8
		x"00",x"01",x"00",x"40",x"00",x"42",x"2C",x"44", -- 0x1AD0
		x"10",x"40",x"40",x"40",x"00",x"02",x"CD",x"00", -- 0x1AD8
		x"02",x"05",x"89",x"10",x"80",x"02",x"58",x"08", -- 0x1AE0
		x"04",x"22",x"00",x"10",x"83",x"0D",x"4A",x"64", -- 0x1AE8
		x"00",x"00",x"80",x"80",x"00",x"80",x"00",x"04", -- 0x1AF0
		x"00",x"80",x"80",x"80",x"00",x"00",x"00",x"00", -- 0x1AF8
		x"40",x"44",x"00",x"05",x"20",x"00",x"04",x"10", -- 0x1B00
		x"10",x"10",x"00",x"40",x"44",x"44",x"00",x"00", -- 0x1B08
		x"82",x"8A",x"00",x"24",x"24",x"84",x"80",x"22", -- 0x1B10
		x"22",x"80",x"10",x"10",x"00",x"04",x"84",x"81", -- 0x1B18
		x"00",x"04",x"44",x"00",x"00",x"01",x"23",x"22", -- 0x1B20
		x"02",x"00",x"10",x"12",x"00",x"00",x"08",x"00", -- 0x1B28
		x"80",x"04",x"04",x"24",x"00",x"00",x"00",x"20", -- 0x1B30
		x"20",x"08",x"00",x"01",x"81",x"80",x"10",x"10", -- 0x1B38
		x"00",x"04",x"44",x"00",x"00",x"01",x"23",x"22", -- 0x1B40
		x"02",x"00",x"10",x"12",x"00",x"00",x"08",x"00", -- 0x1B48
		x"80",x"00",x"04",x"24",x"00",x"00",x"00",x"20", -- 0x1B50
		x"20",x"08",x"00",x"01",x"81",x"80",x"10",x"10", -- 0x1B58
		x"6C",x"D2",x"91",x"11",x"40",x"22",x"08",x"48", -- 0x1B60
		x"44",x"22",x"00",x"11",x"82",x"0C",x"4A",x"64", -- 0x1B68
		x"50",x"A8",x"45",x"D1",x"03",x"04",x"00",x"00", -- 0x1B70
		x"00",x"20",x"24",x"06",x"29",x"4C",x"36",x"0C", -- 0x1B78
		x"81",x"00",x"00",x"02",x"81",x"84",x"02",x"00", -- 0x1B80
		x"02",x"21",x"54",x"21",x"01",x"20",x"60",x"10", -- 0x1B88
		x"00",x"81",x"80",x"40",x"00",x"42",x"2C",x"44", -- 0x1B90
		x"10",x"00",x"42",x"40",x"10",x"1A",x"CD",x"00", -- 0x1B98
		x"01",x"05",x"8C",x"18",x"80",x"02",x"58",x"48", -- 0x1BA0
		x"44",x"22",x"00",x"11",x"82",x"0C",x"4A",x"64", -- 0x1BA8
		x"26",x"A9",x"DD",x"42",x"10",x"0B",x"24",x"00", -- 0x1BB0
		x"04",x"26",x"02",x"02",x"01",x"00",x"80",x"12", -- 0x1BB8
		x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"06", -- 0x1BC0
		x"02",x"05",x"00",x"10",x"08",x"00",x"00",x"00", -- 0x1BC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40", -- 0x1BD0
		x"80",x"40",x"80",x"40",x"20",x"00",x"00",x"00", -- 0x1BD8
		x"00",x"00",x"00",x"00",x"00",x"08",x"04",x"06", -- 0x1BE0
		x"02",x"05",x"00",x"10",x"08",x"00",x"00",x"00", -- 0x1BE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40", -- 0x1BF0
		x"80",x"40",x"80",x"40",x"20",x"00",x"00",x"00", -- 0x1BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"E0", -- 0x1C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"00", -- 0x1C18
		x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"F3", -- 0x1C20
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10", -- 0x1C28
		x"07",x"FF",x"00",x"00",x"FE",x"03",x"00",x"F8", -- 0x1C30
		x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
		x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10", -- 0x1C40
		x"10",x"00",x"00",x"3E",x"41",x"3E",x"00",x"00", -- 0x1C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
		x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- 0x1C58
		x"FF",x"FF",x"FF",x"00",x"00",x"3F",x"FF",x"FF", -- 0x1C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C68
		x"F2",x"C7",x"80",x"00",x"00",x"FF",x"FF",x"FF", -- 0x1C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C78
		x"00",x"00",x"30",x"41",x"A1",x"40",x"20",x"00", -- 0x1C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
		x"50",x"C8",x"90",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
		x"00",x"F8",x"00",x"00",x"80",x"00",x"9E",x"40", -- 0x1CA0
		x"80",x"80",x"80",x"80",x"00",x"00",x"00",x"08", -- 0x1CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
		x"00",x"00",x"83",x"87",x"0F",x"1E",x"1E",x"1E", -- 0x1CB8
		x"2A",x"00",x"02",x"2C",x"2F",x"20",x"3E",x"0F", -- 0x1CC0
		x"07",x"83",x"C1",x"E0",x"70",x"78",x"7C",x"3F", -- 0x1CC8
		x"0E",x"4E",x"8E",x"0E",x"CE",x"0E",x"07",x"07", -- 0x1CD0
		x"07",x"83",x"C1",x"E0",x"F0",x"00",x"00",x"00", -- 0x1CD8
		x"87",x"00",x"00",x"00",x"FF",x"FF",x"02",x"FF", -- 0x1CE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CE8
		x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"FF", -- 0x1CF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"00", -- 0x1D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
		x"00",x"1F",x"20",x"40",x"C2",x"C3",x"C0",x"C0", -- 0x1D20
		x"82",x"20",x"00",x"40",x"20",x"00",x"00",x"00", -- 0x1D28
		x"00",x"FF",x"00",x"00",x"00",x"00",x"20",x"0F", -- 0x1D30
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
		x"00",x"00",x"00",x"00",x"20",x"40",x"00",x"01", -- 0x1D40
		x"00",x"00",x"04",x"00",x"07",x"81",x"C0",x"20", -- 0x1D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
		x"20",x"00",x"80",x"40",x"80",x"00",x"00",x"00", -- 0x1D58
		x"38",x"38",x"38",x"00",x"00",x"00",x"FF",x"FF", -- 0x1D60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D68
		x"FF",x"AB",x"81",x"81",x"00",x"00",x"FF",x"FF", -- 0x1D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D78
		x"0A",x"05",x"0C",x"08",x"10",x"10",x"00",x"00", -- 0x1D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
		x"80",x"00",x"84",x"08",x"08",x"02",x"01",x"03", -- 0x1D90
		x"02",x"04",x"04",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
		x"03",x"0F",x"1F",x"1F",x"3F",x"3C",x"3F",x"38", -- 0x1DA0
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x1DA8
		x"80",x"1F",x"30",x"14",x"0C",x"08",x"FC",x"07", -- 0x1DB0
		x"10",x"1F",x"01",x"01",x"00",x"20",x"3E",x"3F", -- 0x1DB8
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x1DC0
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x1DC8
		x"03",x"03",x"0F",x"03",x"03",x"03",x"03",x"07", -- 0x1DD0
		x"07",x"07",x"07",x"23",x"20",x"00",x"08",x"80", -- 0x1DD8
		x"1F",x"0F",x"0F",x"07",x"07",x"03",x"01",x"FF", -- 0x1DE0
		x"00",x"7D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE8
		x"C3",x"E0",x"F0",x"F8",x"FF",x"FF",x"FF",x"00", -- 0x1DF0
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"00", -- 0x1E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"00", -- 0x1E18
		x"00",x"00",x"1B",x"00",x"24",x"17",x"F7",x"10", -- 0x1E20
		x"07",x"FF",x"F0",x"E0",x"01",x"02",x"02",x"04", -- 0x1E28
		x"00",x"00",x"60",x"08",x"00",x"60",x"68",x"04", -- 0x1E30
		x"F1",x"8F",x"3C",x"F0",x"60",x"41",x"40",x"00", -- 0x1E38
		x"05",x"05",x"05",x"05",x"01",x"01",x"01",x"81", -- 0x1E40
		x"C0",x"F0",x"FC",x"FE",x"00",x"00",x"00",x"00", -- 0x1E48
		x"83",x"00",x"81",x"00",x"80",x"80",x"C0",x"80", -- 0x1E50
		x"00",x"00",x"00",x"3F",x"29",x"29",x"2F",x"31", -- 0x1E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
		x"00",x"00",x"00",x"A0",x"80",x"8A",x"AA",x"20", -- 0x1E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
		x"00",x"00",x"00",x"00",x"22",x"22",x"A4",x"04", -- 0x1E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"94", -- 0x1E80
		x"90",x"55",x"46",x"52",x"58",x"12",x"82",x"81", -- 0x1E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
		x"00",x"20",x"92",x"90",x"91",x"09",x"2B",x"20", -- 0x1E98
		x"00",x"80",x"88",x"A0",x"20",x"20",x"40",x"44", -- 0x1EA0
		x"54",x"18",x"28",x"2A",x"2A",x"82",x"90",x"90", -- 0x1EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"00", -- 0x1EB0
		x"80",x"A0",x"A2",x"50",x"42",x"4A",x"2A",x"28", -- 0x1EB8
		x"80",x"94",x"10",x"50",x"40",x"D4",x"80",x"48", -- 0x1EC0
		x"48",x"0A",x"02",x"33",x"91",x"91",x"88",x"8A", -- 0x1EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08", -- 0x1ED0
		x"00",x"00",x"00",x"00",x"00",x"40",x"40",x"40", -- 0x1ED8
		x"00",x"00",x"00",x"00",x"90",x"80",x"04",x"54", -- 0x1EE0
		x"40",x"A8",x"A4",x"A5",x"20",x"4A",x"6A",x"22", -- 0x1EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80", -- 0x1EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
		x"00",x"00",x"00",x"40",x"40",x"00",x"80",x"90", -- 0x1F08
		x"00",x"00",x"00",x"00",x"40",x"00",x"00",x"00", -- 0x1F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
		x"00",x"00",x"80",x"00",x"20",x"A0",x"40",x"48", -- 0x1F20
		x"10",x"40",x"40",x"A8",x"80",x"10",x"44",x"2A", -- 0x1F28
		x"00",x"00",x"42",x"C4",x"00",x"00",x"00",x"00", -- 0x1F30
		x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00", -- 0x1F38
		x"28",x"40",x"90",x"A2",x"68",x"40",x"14",x"20", -- 0x1F40
		x"48",x"40",x"A0",x"08",x"20",x"80",x"00",x"44", -- 0x1F48
		x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00", -- 0x1F50
		x"00",x"00",x"00",x"00",x"04",x"02",x"00",x"00", -- 0x1F58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
		x"00",x"00",x"00",x"00",x"80",x"80",x"49",x"49", -- 0x1F68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20", -- 0x1F78
		x"29",x"69",x"B2",x"14",x"60",x"8A",x"39",x"A9", -- 0x1F80
		x"C5",x"1F",x"51",x"03",x"2A",x"B5",x"58",x"39", -- 0x1F88
		x"80",x"50",x"00",x"AA",x"A0",x"B1",x"70",x"52", -- 0x1F90
		x"49",x"29",x"A0",x"32",x"50",x"1D",x"54",x"66", -- 0x1F98
		x"66",x"2A",x"B8",x"0A",x"4C",x"05",x"95",x"B2", -- 0x1FA0
		x"4A",x"AE",x"AF",x"A5",x"95",x"D1",x"CA",x"29", -- 0x1FA8
		x"FC",x"3A",x"AD",x"55",x"C1",x"AA",x"F8",x"A3", -- 0x1FB0
		x"95",x"9F",x"51",x"06",x"A8",x"CD",x"96",x"94", -- 0x1FB8
		x"E0",x"00",x"00",x"00",x"80",x"C0",x"00",x"FF", -- 0x1FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC8
		x"25",x"25",x"3E",x"00",x"00",x"00",x"7F",x"FF", -- 0x1FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD8
		x"08",x"10",x"10",x"05",x"02",x"06",x"04",x"08", -- 0x1FE0
		x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FE8
		x"00",x"60",x"80",x"40",x"80",x"40",x"00",x"00", -- 0x1FF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x1FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
