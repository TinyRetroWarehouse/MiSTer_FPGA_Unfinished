-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_M3 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_M3 is


	type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"F3",x"31",x"BE",x"EF",x"C3",x"46",x"01",x"FF", -- 0x0000
		x"E5",x"C5",x"F5",x"C3",x"72",x"01",x"00",x"05", -- 0x0008
		x"E5",x"D5",x"C5",x"F5",x"C3",x"96",x"01",x"70", -- 0x0010
		x"3E",x"02",x"18",x"04",x"70",x"C0",x"3E",x"01", -- 0x0018
		x"F3",x"E5",x"D5",x"C5",x"F5",x"C3",x"FC",x"00", -- 0x0020
		x"F3",x"E5",x"D5",x"C5",x"F5",x"C3",x"F3",x"00", -- 0x0028
		x"F3",x"CD",x"39",x"01",x"72",x"C3",x"82",x"00", -- 0x0030
		x"F3",x"E5",x"D5",x"C5",x"F5",x"CD",x"3C",x"01", -- 0x0038
		x"36",x"40",x"23",x"72",x"23",x"71",x"23",x"70", -- 0x0040
		x"C3",x"CD",x"00",x"21",x"C0",x"EF",x"01",x"00", -- 0x0048
		x"10",x"11",x"04",x"00",x"AF",x"CB",x"4E",x"28", -- 0x0050
		x"0B",x"23",x"35",x"2B",x"20",x"06",x"36",x"30", -- 0x0058
		x"B9",x"20",x"01",x"48",x"19",x"10",x"EE",x"B9", -- 0x0060
		x"CA",x"CD",x"00",x"3A",x"BF",x"EF",x"47",x"CD", -- 0x0068
		x"3C",x"01",x"7E",x"FE",x"20",x"C2",x"84",x"00", -- 0x0070
		x"3E",x"10",x"91",x"B8",x"DA",x"2E",x"01",x"C3", -- 0x0078
		x"CD",x"00",x"23",x"72",x"31",x"BE",x"EF",x"FB", -- 0x0080
		x"21",x"C0",x"EF",x"01",x"00",x"10",x"11",x"04", -- 0x0088
		x"00",x"7E",x"FE",x"20",x"30",x"06",x"0C",x"19", -- 0x0090
		x"10",x"F7",x"18",x"EB",x"F3",x"79",x"32",x"BF", -- 0x0098
		x"EF",x"7E",x"36",x"20",x"23",x"72",x"23",x"5E", -- 0x00A0
		x"23",x"56",x"FE",x"40",x"38",x"13",x"7D",x"E6", -- 0x00A8
		x"3C",x"0F",x"4F",x"06",x"00",x"21",x"D3",x"00", -- 0x00B0
		x"09",x"7E",x"23",x"66",x"6F",x"F9",x"EB",x"FB", -- 0x00B8
		x"E9",x"EB",x"F9",x"F1",x"C1",x"D1",x"E1",x"FD", -- 0x00C0
		x"E1",x"DD",x"E1",x"D9",x"08",x"F1",x"C1",x"D1", -- 0x00C8
		x"E1",x"FB",x"C9",x"98",x"EF",x"68",x"EF",x"38", -- 0x00D0
		x"EF",x"08",x"EF",x"D8",x"EE",x"A8",x"EE",x"78", -- 0x00D8
		x"EE",x"48",x"EE",x"18",x"EE",x"E8",x"ED",x"B8", -- 0x00E0
		x"ED",x"88",x"ED",x"58",x"ED",x"28",x"ED",x"F8", -- 0x00E8
		x"EC",x"C8",x"EC",x"CD",x"3C",x"01",x"72",x"23", -- 0x00F0
		x"72",x"C3",x"CD",x"00",x"CD",x"39",x"01",x"36", -- 0x00F8
		x"12",x"23",x"70",x"2B",x"AF",x"08",x"23",x"23", -- 0x0100
		x"EB",x"21",x"F4",x"FF",x"39",x"EB",x"73",x"23", -- 0x0108
		x"72",x"D9",x"DD",x"E5",x"FD",x"E5",x"E5",x"D5", -- 0x0110
		x"C5",x"F5",x"08",x"CA",x"84",x"00",x"CD",x"39", -- 0x0118
		x"01",x"C3",x"A1",x"00",x"3A",x"BF",x"EF",x"47", -- 0x0120
		x"F1",x"F5",x"B8",x"D2",x"CD",x"00",x"32",x"BF", -- 0x0128
		x"EF",x"78",x"CD",x"3C",x"01",x"3C",x"C3",x"05", -- 0x0130
		x"01",x"3A",x"BF",x"EF",x"21",x"C0",x"EF",x"07", -- 0x0138
		x"07",x"5F",x"AF",x"57",x"19",x"C9",x"CD",x"A7", -- 0x0140
		x"02",x"21",x"00",x"E0",x"01",x"00",x"10",x"36", -- 0x0148
		x"00",x"23",x"0B",x"78",x"B1",x"20",x"F8",x"CD", -- 0x0150
		x"16",x"04",x"3A",x"04",x"C0",x"CB",x"5F",x"20", -- 0x0158
		x"08",x"3E",x"02",x"32",x"06",x"C8",x"C3",x"FE", -- 0x0160
		x"AC",x"01",x"B5",x"02",x"3E",x"06",x"FF",x"C3", -- 0x0168
		x"84",x"00",x"3A",x"04",x"C0",x"07",x"30",x"FA", -- 0x0170
		x"2A",x"20",x"E2",x"7E",x"0E",x"FF",x"3C",x"28", -- 0x0178
		x"09",x"3D",x"4F",x"36",x"FF",x"23",x"7D",x"E6", -- 0x0180
		x"1F",x"6F",x"22",x"20",x"E2",x"79",x"32",x"00", -- 0x0188
		x"C8",x"F1",x"C1",x"E1",x"FB",x"C9",x"21",x"00", -- 0x0190
		x"EB",x"11",x"00",x"CC",x"01",x"80",x"00",x"ED", -- 0x0198
		x"B0",x"3A",x"C7",x"EB",x"CB",x"47",x"28",x"33", -- 0x01A0
		x"EE",x"02",x"32",x"C7",x"EB",x"E6",x"02",x"28", -- 0x01A8
		x"2A",x"2A",x"D2",x"E0",x"23",x"22",x"D2",x"E0", -- 0x01B0
		x"22",x"02",x"C8",x"7D",x"E6",x"7F",x"7D",x"20", -- 0x01B8
		x"05",x"21",x"A4",x"E9",x"36",x"01",x"E6",x"0F", -- 0x01C0
		x"C2",x"DB",x"01",x"21",x"DF",x"EB",x"CB",x"C6", -- 0x01C8
		x"23",x"23",x"ED",x"5B",x"C2",x"EB",x"01",x"1E", -- 0x01D0
		x"00",x"ED",x"B0",x"3E",x"02",x"C3",x"4B",x"00", -- 0x01D8
		x"16",x"30",x"72",x"23",x"0B",x"79",x"B0",x"20", -- 0x01E0
		x"F9",x"C9",x"06",x"01",x"18",x"01",x"1A",x"77", -- 0x01E8
		x"13",x"C5",x"01",x"20",x"00",x"09",x"C1",x"10", -- 0x01F0
		x"F5",x"C9",x"0E",x"00",x"1A",x"81",x"0E",x"00", -- 0x01F8
		x"86",x"FE",x"0A",x"38",x"03",x"0C",x"D6",x"0A", -- 0x0200
		x"12",x"1B",x"2B",x"10",x"EF",x"C9",x"0E",x"00", -- 0x0208
		x"7E",x"81",x"4F",x"1A",x"91",x"0E",x"00",x"30", -- 0x0210
		x"03",x"0C",x"C6",x"0A",x"12",x"1B",x"2B",x"10", -- 0x0218
		x"EF",x"C9",x"46",x"23",x"4E",x"AF",x"B9",x"C8", -- 0x0220
		x"23",x"5E",x"23",x"56",x"23",x"EB",x"B8",x"20", -- 0x0228
		x"08",x"C5",x"41",x"CD",x"EE",x"01",x"C1",x"18", -- 0x0230
		x"0B",x"C5",x"DF",x"06",x"01",x"CD",x"EE",x"01", -- 0x0238
		x"C1",x"0D",x"20",x"F5",x"EB",x"18",x"DD",x"0E", -- 0x0240
		x"30",x"C5",x"71",x"01",x"20",x"00",x"09",x"C1", -- 0x0248
		x"10",x"F7",x"C9",x"C5",x"E5",x"72",x"23",x"0D", -- 0x0250
		x"20",x"FB",x"E1",x"01",x"20",x"00",x"09",x"C1", -- 0x0258
		x"10",x"F1",x"C9",x"05",x"1A",x"B7",x"20",x"09", -- 0x0260
		x"C5",x"3E",x"30",x"CD",x"EA",x"01",x"C1",x"10", -- 0x0268
		x"F3",x"04",x"C3",x"EE",x"01",x"EB",x"C5",x"D5", -- 0x0270
		x"06",x"00",x"ED",x"B0",x"EB",x"0E",x"20",x"E1", -- 0x0278
		x"09",x"C1",x"10",x"F1",x"C9",x"AF",x"6F",x"67", -- 0x0280
		x"22",x"D0",x"E0",x"22",x"D2",x"E0",x"32",x"D5", -- 0x0288
		x"E0",x"22",x"00",x"C8",x"22",x"02",x"C8",x"32", -- 0x0290
		x"05",x"C8",x"C9",x"AF",x"32",x"D5",x"E0",x"32", -- 0x0298
		x"05",x"C8",x"C9",x"3E",x"07",x"18",x"F5",x"21", -- 0x02A0
		x"00",x"EB",x"11",x"01",x"EB",x"01",x"7F",x"00", -- 0x02A8
		x"36",x"00",x"ED",x"B0",x"C9",x"21",x"00",x"00", -- 0x02B0
		x"22",x"18",x"E0",x"22",x"1A",x"E0",x"22",x"16", -- 0x02B8
		x"E0",x"3E",x"1E",x"32",x"C0",x"E9",x"CD",x"A7", -- 0x02C0
		x"02",x"CD",x"B6",x"11",x"CD",x"16",x"04",x"CD", -- 0x02C8
		x"E0",x"11",x"3E",x"10",x"32",x"D4",x"E0",x"CD", -- 0x02D0
		x"8D",x"11",x"CD",x"FD",x"2C",x"CD",x"C7",x"03", -- 0x02D8
		x"DD",x"21",x"2A",x"04",x"CD",x"19",x"2D",x"21", -- 0x02E0
		x"18",x"E0",x"01",x"03",x"C0",x"16",x"80",x"CD", -- 0x02E8
		x"16",x"03",x"21",x"1A",x"E0",x"01",x"04",x"C0", -- 0x02F0
		x"16",x"40",x"CD",x"16",x"03",x"CD",x"A2",x"03", -- 0x02F8
		x"21",x"0C",x"E0",x"34",x"20",x"0A",x"23",x"34", -- 0x0300
		x"20",x"06",x"23",x"34",x"20",x"02",x"23",x"34", -- 0x0308
		x"06",x"01",x"DF",x"C3",x"E7",x"02",x"0A",x"E6", -- 0x0310
		x"07",x"20",x"08",x"21",x"00",x"02",x"22",x"10", -- 0x0318
		x"E0",x"18",x"5C",x"7E",x"B7",x"3A",x"00",x"C0", -- 0x0320
		x"20",x"04",x"A2",x"C0",x"18",x"06",x"A2",x"7E", -- 0x0328
		x"20",x"04",x"3C",x"C8",x"34",x"C9",x"36",x"00", -- 0x0330
		x"FE",x"19",x"D0",x"D9",x"21",x"20",x"E0",x"34", -- 0x0338
		x"D9",x"23",x"34",x"CB",x"41",x"11",x"9D",x"78", -- 0x0340
		x"20",x"03",x"11",x"AD",x"78",x"0A",x"E6",x"07", -- 0x0348
		x"07",x"4F",x"06",x"00",x"EB",x"09",x"4E",x"23", -- 0x0350
		x"46",x"1A",x"B9",x"D8",x"3A",x"10",x"E0",x"FE", -- 0x0358
		x"09",x"38",x"07",x"3A",x"11",x"E0",x"80",x"FE", -- 0x0360
		x"0A",x"D0",x"60",x"AF",x"6F",x"22",x"12",x"E0", -- 0x0368
		x"2B",x"1A",x"91",x"12",x"21",x"13",x"E0",x"11", -- 0x0370
		x"11",x"E0",x"06",x"02",x"CD",x"FA",x"01",x"3A", -- 0x0378
		x"00",x"E0",x"0F",x"D4",x"0C",x"12",x"21",x"00", -- 0x0380
		x"E0",x"7E",x"07",x"38",x"08",x"36",x"80",x"3E", -- 0x0388
		x"00",x"01",x"46",x"13",x"FF",x"CB",x"4E",x"C0", -- 0x0390
		x"3E",x"38",x"32",x"15",x"E0",x"0E",x"0A",x"C3", -- 0x0398
		x"78",x"11",x"21",x"16",x"E0",x"16",x"10",x"7E", -- 0x03A0
		x"B7",x"3A",x"00",x"C0",x"20",x"04",x"A2",x"C0", -- 0x03A8
		x"18",x"06",x"A2",x"7E",x"20",x"04",x"3C",x"C8", -- 0x03B0
		x"34",x"C9",x"36",x"00",x"11",x"17",x"E0",x"3E", -- 0x03B8
		x"01",x"12",x"01",x"01",x"01",x"18",x"95",x"AF", -- 0x03C0
		x"0E",x"25",x"21",x"00",x"E8",x"77",x"3C",x"23", -- 0x03C8
		x"36",x"00",x"23",x"36",x"00",x"23",x"71",x"23", -- 0x03D0
		x"36",x"00",x"23",x"08",x"79",x"E6",x"0F",x"20", -- 0x03D8
		x"06",x"79",x"D6",x"10",x"F6",x"0A",x"4F",x"0D", -- 0x03E0
		x"06",x"08",x"36",x"30",x"23",x"10",x"FB",x"06", -- 0x03E8
		x"03",x"36",x"00",x"23",x"10",x"FB",x"08",x"FE", -- 0x03F0
		x"19",x"38",x"D2",x"11",x"01",x"E8",x"21",x"CE", -- 0x03F8
		x"A3",x"3E",x"0A",x"01",x"0C",x"00",x"ED",x"B0", -- 0x0400
		x"13",x"13",x"13",x"13",x"3D",x"20",x"F4",x"21", -- 0x0408
		x"00",x"04",x"22",x"42",x"E0",x"C9",x"21",x"00", -- 0x0410
		x"E2",x"22",x"22",x"E2",x"22",x"20",x"E2",x"11", -- 0x0418
		x"01",x"E2",x"36",x"FF",x"01",x"1F",x"00",x"ED", -- 0x0420
		x"B0",x"C9",x"03",x"6F",x"0F",x"00",x"40",x"0F", -- 0x0428
		x"0A",x"12",x"71",x"0F",x"3A",x"43",x"E1",x"B7", -- 0x0430
		x"C2",x"69",x"05",x"3A",x"76",x"E1",x"B7",x"C2", -- 0x0438
		x"37",x"05",x"21",x"54",x"E1",x"35",x"C2",x"46", -- 0x0440
		x"05",x"36",x"01",x"EB",x"3A",x"70",x"E1",x"21", -- 0x0448
		x"71",x"E1",x"BE",x"D2",x"46",x"05",x"3A",x"1B", -- 0x0450
		x"E1",x"B7",x"C2",x"78",x"08",x"3A",x"45",x"E1", -- 0x0458
		x"B7",x"CA",x"46",x"05",x"47",x"3A",x"53",x"E1", -- 0x0460
		x"12",x"3A",x"EF",x"E0",x"3C",x"32",x"EF",x"E0", -- 0x0468
		x"0F",x"E6",x"0F",x"B8",x"38",x"03",x"90",x"18", -- 0x0470
		x"FA",x"07",x"5F",x"16",x"00",x"21",x"00",x"E7", -- 0x0478
		x"19",x"7E",x"FE",x"FF",x"CA",x"2E",x"05",x"07", -- 0x0480
		x"DA",x"24",x"05",x"11",x"48",x"E1",x"C5",x"01", -- 0x0488
		x"02",x"00",x"F3",x"ED",x"B0",x"FB",x"C1",x"CD", -- 0x0490
		x"8D",x"0C",x"DA",x"69",x"05",x"16",x"03",x"CD", -- 0x0498
		x"51",x"0C",x"38",x"7A",x"CD",x"A8",x"0C",x"ED", -- 0x04A0
		x"5B",x"48",x"E1",x"7B",x"E6",x"03",x"4F",x"0F", -- 0x04A8
		x"0F",x"FD",x"77",x"01",x"21",x"70",x"E1",x"79", -- 0x04B0
		x"0F",x"30",x"14",x"7A",x"FD",x"77",x"05",x"FD", -- 0x04B8
		x"36",x"21",x"01",x"3A",x"03",x"E1",x"FE",x"10", -- 0x04C0
		x"3E",x"00",x"38",x"28",x"3C",x"18",x"25",x"0F", -- 0x04C8
		x"30",x"05",x"7A",x"E6",x"01",x"18",x"1D",x"7A", -- 0x04D0
		x"FD",x"77",x"05",x"FE",x"18",x"3E",x"01",x"30", -- 0x04D8
		x"0A",x"3A",x"03",x"E1",x"FE",x"07",x"3E",x"01", -- 0x04E0
		x"30",x"01",x"AF",x"FD",x"77",x"21",x"7B",x"07", -- 0x04E8
		x"07",x"07",x"E6",x"03",x"34",x"FD",x"77",x"1D", -- 0x04F0
		x"FD",x"77",x"1A",x"07",x"FD",x"77",x"0D",x"AF", -- 0x04F8
		x"FD",x"77",x"03",x"FD",x"77",x"08",x"FD",x"36", -- 0x0500
		x"00",x"01",x"7E",x"21",x"71",x"E1",x"BE",x"38", -- 0x0508
		x"35",x"2A",x"72",x"E1",x"22",x"74",x"E1",x"3E", -- 0x0510
		x"01",x"32",x"76",x"E1",x"18",x"28",x"FD",x"36", -- 0x0518
		x"00",x"00",x"18",x"45",x"11",x"02",x"00",x"19", -- 0x0520
		x"7D",x"FE",x"20",x"DA",x"31",x"05",x"21",x"00", -- 0x0528
		x"E7",x"05",x"C2",x"81",x"04",x"18",x"0F",x"2A", -- 0x0530
		x"74",x"E1",x"2B",x"22",x"74",x"E1",x"7D",x"B4", -- 0x0538
		x"20",x"04",x"AF",x"32",x"76",x"E1",x"3A",x"E0", -- 0x0540
		x"E7",x"B7",x"C4",x"6F",x"05",x"3A",x"B0",x"E7", -- 0x0548
		x"B7",x"C4",x"BC",x"0B",x"3A",x"00",x"EC",x"B7", -- 0x0550
		x"C4",x"2A",x"0B",x"3A",x"07",x"E1",x"B7",x"C4", -- 0x0558
		x"01",x"0B",x"3A",x"14",x"E1",x"B7",x"C4",x"B9", -- 0x0560
		x"08",x"06",x"02",x"DF",x"C3",x"34",x"04",x"3A", -- 0x0568
		x"E0",x"E7",x"E6",x"40",x"C2",x"B1",x"05",x"3A", -- 0x0570
		x"E1",x"E7",x"E6",x"E0",x"FE",x"60",x"3E",x"05", -- 0x0578
		x"20",x"02",x"3E",x"0A",x"32",x"ED",x"E7",x"3A", -- 0x0580
		x"E2",x"E7",x"4F",x"3A",x"ED",x"E7",x"91",x"28", -- 0x0588
		x"1B",x"47",x"C5",x"CD",x"8D",x"0C",x"C1",x"D8", -- 0x0590
		x"CD",x"5D",x"07",x"CD",x"9B",x"07",x"3A",x"ED", -- 0x0598
		x"E7",x"4F",x"3A",x"E2",x"E7",x"3C",x"32",x"E2", -- 0x05A0
		x"E7",x"B9",x"38",x"05",x"21",x"E0",x"E7",x"CB", -- 0x05A8
		x"F6",x"3A",x"E0",x"E7",x"E6",x"20",x"C2",x"36", -- 0x05B0
		x"06",x"32",x"E4",x"E7",x"3A",x"ED",x"E7",x"47", -- 0x05B8
		x"21",x"C0",x"E7",x"CB",x"46",x"23",x"CA",x"CE", -- 0x05C0
		x"05",x"CB",x"7E",x"C2",x"DB",x"05",x"3A",x"E4", -- 0x05C8
		x"E7",x"3C",x"32",x"E4",x"E7",x"23",x"10",x"EB", -- 0x05D0
		x"C3",x"29",x"06",x"E5",x"C5",x"01",x"13",x"06", -- 0x05D8
		x"21",x"F9",x"05",x"3A",x"E1",x"E7",x"E6",x"E0", -- 0x05E0
		x"FE",x"60",x"20",x"03",x"21",x"03",x"06",x"C5", -- 0x05E8
		x"3A",x"E0",x"E7",x"E6",x"0F",x"CD",x"36",x"19", -- 0x05F0
		x"E9",x"AA",x"07",x"C2",x"07",x"E1",x"07",x"E1", -- 0x05F8
		x"07",x"02",x"08",x"43",x"08",x"54",x"08",x"5F", -- 0x0600
		x"08",x"54",x"08",x"63",x"08",x"67",x"08",x"5F", -- 0x0608
		x"08",x"3F",x"08",x"16",x"03",x"CD",x"51",x"0C", -- 0x0610
		x"C1",x"3E",x"80",x"38",x"0A",x"3A",x"E3",x"E7", -- 0x0618
		x"3C",x"32",x"E3",x"E7",x"7D",x"E6",x"1F",x"E1", -- 0x0620
		x"77",x"21",x"ED",x"E7",x"3A",x"E3",x"E7",x"BE", -- 0x0628
		x"D8",x"21",x"E0",x"E7",x"CB",x"EE",x"3A",x"E0", -- 0x0630
		x"E7",x"57",x"2F",x"E6",x"60",x"C0",x"AF",x"32", -- 0x0638
		x"E4",x"E7",x"CD",x"67",x"07",x"23",x"7E",x"CD", -- 0x0640
		x"32",x"5F",x"DD",x"77",x"0B",x"2A",x"E0",x"E7", -- 0x0648
		x"7D",x"E6",x"0F",x"DD",x"77",x"02",x"DD",x"74", -- 0x0650
		x"08",x"21",x"D1",x"7F",x"3A",x"E1",x"E7",x"E6", -- 0x0658
		x"E0",x"FE",x"60",x"20",x"03",x"21",x"B4",x"AA", -- 0x0660
		x"3A",x"E0",x"E7",x"E6",x"0F",x"07",x"4F",x"06", -- 0x0668
		x"00",x"09",x"7E",x"23",x"66",x"6F",x"3A",x"E1", -- 0x0670
		x"E7",x"E6",x"E0",x"FE",x"60",x"28",x"0A",x"3A", -- 0x0678
		x"E4",x"E7",x"07",x"4F",x"09",x"7E",x"23",x"66", -- 0x0680
		x"6F",x"7E",x"DD",x"77",x"16",x"23",x"7E",x"DD", -- 0x0688
		x"77",x"19",x"23",x"DD",x"75",x"10",x"DD",x"74", -- 0x0690
		x"11",x"DD",x"36",x"1A",x"02",x"DD",x"36",x"1D", -- 0x0698
		x"02",x"2A",x"E8",x"E7",x"DD",x"75",x"1E",x"DD", -- 0x06A0
		x"74",x"1F",x"21",x"F2",x"86",x"3A",x"E1",x"E7", -- 0x06A8
		x"E6",x"E0",x"FE",x"60",x"20",x"03",x"21",x"3E", -- 0x06B0
		x"B0",x"CD",x"83",x"07",x"3A",x"E6",x"E7",x"86", -- 0x06B8
		x"DD",x"77",x"0F",x"23",x"3A",x"E5",x"E7",x"86", -- 0x06C0
		x"DD",x"77",x"0E",x"23",x"3A",x"E7",x"E7",x"DD", -- 0x06C8
		x"77",x"13",x"7E",x"E6",x"7F",x"DD",x"77",x"14", -- 0x06D0
		x"7E",x"E6",x"80",x"0F",x"0F",x"DD",x"B6",x"02", -- 0x06D8
		x"DD",x"77",x"02",x"23",x"7E",x"DD",x"77",x"0D", -- 0x06E0
		x"DD",x"7E",x"19",x"CD",x"E6",x"32",x"CD",x"0A", -- 0x06E8
		x"42",x"DD",x"77",x"0C",x"AF",x"DD",x"77",x"03", -- 0x06F0
		x"DD",x"77",x"0A",x"DD",x"77",x"01",x"DD",x"36", -- 0x06F8
		x"04",x"01",x"DD",x"7E",x"08",x"E6",x"F0",x"21", -- 0x0700
		x"E4",x"E7",x"B6",x"DD",x"77",x"08",x"34",x"7E", -- 0x0708
		x"21",x"ED",x"E7",x"BE",x"DA",x"42",x"06",x"AF", -- 0x0710
		x"32",x"E0",x"E7",x"32",x"E2",x"E7",x"32",x"E3", -- 0x0718
		x"E7",x"32",x"E4",x"E7",x"2A",x"E8",x"E7",x"3A", -- 0x0720
		x"ED",x"E7",x"77",x"23",x"77",x"23",x"7D",x"E6", -- 0x0728
		x"0F",x"20",x"03",x"21",x"F0",x"E7",x"22",x"E8", -- 0x0730
		x"E7",x"CD",x"67",x"07",x"DD",x"36",x"00",x"11", -- 0x0738
		x"3A",x"E4",x"E7",x"3C",x"32",x"E4",x"E7",x"21", -- 0x0740
		x"ED",x"E7",x"BE",x"38",x"EC",x"21",x"C0",x"E7", -- 0x0748
		x"3E",x"0A",x"11",x"00",x"80",x"47",x"73",x"23", -- 0x0750
		x"72",x"23",x"10",x"FA",x"C9",x"21",x"C0",x"E7", -- 0x0758
		x"59",x"CB",x"03",x"16",x"00",x"19",x"C9",x"21", -- 0x0760
		x"C0",x"E7",x"3A",x"E4",x"E7",x"07",x"4F",x"06", -- 0x0768
		x"00",x"09",x"7E",x"E6",x"FC",x"87",x"CB",x"10", -- 0x0770
		x"87",x"CB",x"10",x"4F",x"DD",x"21",x"00",x"E4", -- 0x0778
		x"DD",x"09",x"C9",x"3A",x"E4",x"E7",x"57",x"3A", -- 0x0780
		x"E0",x"E7",x"E6",x"0F",x"07",x"4F",x"06",x"00", -- 0x0788
		x"09",x"7E",x"23",x"66",x"6F",x"7A",x"07",x"07", -- 0x0790
		x"4F",x"09",x"C9",x"FD",x"E5",x"D1",x"7B",x"CB", -- 0x0798
		x"0A",x"1F",x"CB",x"0A",x"1F",x"E6",x"FC",x"3C", -- 0x07A0
		x"77",x"C9",x"3A",x"E0",x"E7",x"E6",x"10",x"C0", -- 0x07A8
		x"3A",x"0C",x"E0",x"E6",x"0F",x"C6",x"D0",x"32", -- 0x07B0
		x"E6",x"E7",x"3E",x"10",x"32",x"E7",x"E7",x"C3", -- 0x07B8
		x"D7",x"07",x"3A",x"E0",x"E7",x"E6",x"10",x"C0", -- 0x07C0
		x"3A",x"0C",x"E0",x"E6",x"1F",x"C6",x"C0",x"32", -- 0x07C8
		x"E6",x"E7",x"3E",x"08",x"32",x"E7",x"E7",x"AF", -- 0x07D0
		x"32",x"E5",x"E7",x"21",x"E0",x"E7",x"CB",x"E6", -- 0x07D8
		x"C9",x"3A",x"E0",x"E7",x"E6",x"10",x"C0",x"2A", -- 0x07E0
		x"EC",x"E0",x"23",x"24",x"22",x"EC",x"E0",x"7D", -- 0x07E8
		x"E6",x"1F",x"C6",x"80",x"32",x"E6",x"E7",x"7C", -- 0x07F0
		x"E6",x"0F",x"C6",x"08",x"32",x"E7",x"E7",x"C3", -- 0x07F8
		x"D7",x"07",x"3A",x"E0",x"E7",x"E6",x"10",x"C0", -- 0x0800
		x"2A",x"E8",x"E0",x"23",x"24",x"22",x"E8",x"E0", -- 0x0808
		x"01",x"38",x"5C",x"3A",x"0E",x"E1",x"FE",x"3C", -- 0x0810
		x"38",x"0D",x"FE",x"94",x"30",x"09",x"01",x"1C", -- 0x0818
		x"78",x"FE",x"46",x"38",x"02",x"06",x"5C",x"7D", -- 0x0820
		x"A1",x"80",x"32",x"E5",x"E7",x"7C",x"E6",x"0F", -- 0x0828
		x"C6",x"08",x"32",x"E7",x"E7",x"AF",x"32",x"E6", -- 0x0830
		x"E7",x"21",x"E0",x"E7",x"CB",x"E6",x"C9",x"3E", -- 0x0838
		x"E0",x"18",x"02",x"3E",x"48",x"32",x"E6",x"E7", -- 0x0840
		x"AF",x"32",x"E5",x"E7",x"3E",x"08",x"32",x"E7", -- 0x0848
		x"E7",x"C3",x"39",x"08",x"3E",x"18",x"32",x"E5", -- 0x0850
		x"E7",x"AF",x"32",x"E6",x"E7",x"18",x"ED",x"3E", -- 0x0858
		x"28",x"18",x"F3",x"3E",x"A0",x"18",x"DE",x"3E", -- 0x0860
		x"18",x"32",x"E5",x"E7",x"3E",x"F0",x"32",x"E6", -- 0x0868
		x"E7",x"3E",x"10",x"32",x"E7",x"E7",x"18",x"D4", -- 0x0870
		x"CD",x"8D",x"0C",x"DA",x"69",x"05",x"16",x"03", -- 0x0878
		x"CD",x"51",x"0C",x"38",x"2D",x"CD",x"A8",x"0C", -- 0x0880
		x"3A",x"53",x"E1",x"32",x"54",x"E1",x"21",x"1B", -- 0x0888
		x"E1",x"35",x"AF",x"FD",x"77",x"1A",x"FD",x"77", -- 0x0890
		x"1D",x"FD",x"77",x"0D",x"FD",x"36",x"01",x"20", -- 0x0898
		x"FD",x"77",x"03",x"FD",x"77",x"08",x"FD",x"36", -- 0x08A0
		x"00",x"01",x"21",x"70",x"E1",x"34",x"7E",x"C3", -- 0x08A8
		x"0B",x"05",x"FD",x"36",x"00",x"00",x"C3",x"69", -- 0x08B0
		x"05",x"3A",x"14",x"E1",x"CB",x"57",x"C2",x"07", -- 0x08B8
		x"09",x"3A",x"15",x"E1",x"4F",x"CB",x"7F",x"20", -- 0x08C0
		x"05",x"79",x"E6",x"07",x"18",x"0B",x"07",x"07", -- 0x08C8
		x"07",x"E6",x"03",x"FE",x"03",x"20",x"01",x"3C", -- 0x08D0
		x"3C",x"32",x"4E",x"EC",x"3A",x"48",x"EC",x"4F", -- 0x08D8
		x"3A",x"4E",x"EC",x"91",x"28",x"1C",x"47",x"C5", -- 0x08E0
		x"CD",x"8D",x"0C",x"C1",x"D8",x"21",x"30",x"EC", -- 0x08E8
		x"CD",x"60",x"07",x"CD",x"9B",x"07",x"21",x"4E", -- 0x08F0
		x"EC",x"3A",x"48",x"EC",x"3C",x"32",x"48",x"EC", -- 0x08F8
		x"BE",x"D8",x"21",x"14",x"E1",x"CB",x"D6",x"3A", -- 0x0900
		x"14",x"E1",x"E6",x"02",x"C2",x"79",x"09",x"32", -- 0x0908
		x"4A",x"EC",x"3A",x"4E",x"EC",x"47",x"21",x"30", -- 0x0910
		x"EC",x"DD",x"21",x"3E",x"EC",x"CB",x"46",x"23", -- 0x0918
		x"CA",x"2F",x"09",x"CB",x"7E",x"C2",x"41",x"09", -- 0x0920
		x"DD",x"CB",x"00",x"7E",x"C2",x"3E",x"09",x"3A", -- 0x0928
		x"4A",x"EC",x"3C",x"32",x"4A",x"EC",x"DD",x"23", -- 0x0930
		x"23",x"10",x"E2",x"C3",x"68",x"09",x"DD",x"E5", -- 0x0938
		x"E1",x"E5",x"C5",x"21",x"54",x"09",x"E5",x"3A", -- 0x0940
		x"15",x"E1",x"E6",x"80",x"07",x"CD",x"F7",x"66", -- 0x0948
		x"7A",x"0A",x"A5",x"0A",x"CD",x"51",x"0C",x"C1", -- 0x0950
		x"3E",x"80",x"38",x"0A",x"3A",x"49",x"EC",x"3C", -- 0x0958
		x"32",x"49",x"EC",x"7D",x"E6",x"1F",x"E1",x"77", -- 0x0960
		x"3A",x"4E",x"EC",x"E6",x"07",x"07",x"57",x"3A", -- 0x0968
		x"49",x"EC",x"BA",x"D8",x"21",x"14",x"E1",x"CB", -- 0x0970
		x"CE",x"3A",x"14",x"E1",x"57",x"2F",x"E6",x"06", -- 0x0978
		x"C0",x"AF",x"32",x"4A",x"EC",x"21",x"30",x"EC", -- 0x0980
		x"3A",x"4A",x"EC",x"CD",x"6D",x"07",x"23",x"7E", -- 0x0988
		x"CD",x"32",x"5F",x"DD",x"77",x"0B",x"3A",x"4A", -- 0x0990
		x"EC",x"4F",x"06",x"00",x"21",x"3E",x"EC",x"09", -- 0x0998
		x"7E",x"CD",x"32",x"5F",x"DD",x"77",x"2B",x"3A", -- 0x09A0
		x"15",x"E1",x"E6",x"98",x"DD",x"77",x"08",x"3A", -- 0x09A8
		x"14",x"E1",x"E6",x"60",x"07",x"07",x"07",x"DD", -- 0x09B0
		x"77",x"1A",x"DD",x"77",x"1D",x"CD",x"51",x"0A", -- 0x09B8
		x"3A",x"4C",x"EC",x"86",x"DD",x"77",x"0F",x"23", -- 0x09C0
		x"3A",x"4B",x"EC",x"86",x"DD",x"77",x"0E",x"23", -- 0x09C8
		x"3A",x"4D",x"EC",x"DD",x"77",x"13",x"7E",x"E6", -- 0x09D0
		x"3F",x"07",x"07",x"DD",x"77",x"14",x"7E",x"E6", -- 0x09D8
		x"80",x"0F",x"0F",x"4F",x"3A",x"15",x"E1",x"E6", -- 0x09E0
		x"07",x"B1",x"DD",x"77",x"02",x"23",x"DD",x"7E", -- 0x09E8
		x"1D",x"07",x"B6",x"DD",x"77",x"0D",x"AF",x"DD", -- 0x09F0
		x"77",x"03",x"DD",x"77",x"0A",x"DD",x"36",x"01", -- 0x09F8
		x"C0",x"DD",x"36",x"04",x"01",x"21",x"4A",x"EC", -- 0x0A00
		x"DD",x"7E",x"08",x"B6",x"DD",x"77",x"08",x"34", -- 0x0A08
		x"7E",x"21",x"4E",x"EC",x"BE",x"DA",x"85",x"09", -- 0x0A10
		x"AF",x"32",x"14",x"E1",x"32",x"48",x"EC",x"32", -- 0x0A18
		x"49",x"EC",x"32",x"4A",x"EC",x"21",x"30",x"EC", -- 0x0A20
		x"3A",x"4A",x"EC",x"CD",x"6D",x"07",x"DD",x"36", -- 0x0A28
		x"00",x"11",x"3A",x"4A",x"EC",x"3C",x"32",x"4A", -- 0x0A30
		x"EC",x"21",x"4E",x"EC",x"BE",x"38",x"E6",x"21", -- 0x0A38
		x"30",x"EC",x"3E",x"07",x"CD",x"52",x"07",x"06", -- 0x0A40
		x"07",x"21",x"3E",x"EC",x"72",x"23",x"10",x"FC", -- 0x0A48
		x"C9",x"3A",x"4A",x"EC",x"57",x"3A",x"15",x"E1", -- 0x0A50
		x"5F",x"CB",x"7F",x"28",x"08",x"21",x"6B",x"B2", -- 0x0A58
		x"E6",x"07",x"C3",x"8A",x"07",x"21",x"1B",x"B3", -- 0x0A60
		x"3A",x"4B",x"EC",x"FE",x"80",x"38",x"03",x"21", -- 0x0A68
		x"2F",x"B3",x"7A",x"07",x"07",x"4F",x"06",x"00", -- 0x0A70
		x"09",x"C9",x"16",x"03",x"3A",x"14",x"E1",x"E6", -- 0x0A78
		x"08",x"C0",x"3A",x"45",x"EC",x"3C",x"32",x"45", -- 0x0A80
		x"EC",x"0F",x"06",x"20",x"38",x"02",x"06",x"B0", -- 0x0A88
		x"E6",x"0F",x"80",x"32",x"4B",x"EC",x"AF",x"32", -- 0x0A90
		x"4C",x"EC",x"3E",x"10",x"32",x"4D",x"EC",x"21", -- 0x0A98
		x"14",x"E1",x"CB",x"DE",x"C9",x"16",x"03",x"3A", -- 0x0AA0
		x"14",x"E1",x"E6",x"08",x"C0",x"3A",x"15",x"E1", -- 0x0AA8
		x"E6",x"07",x"FE",x"04",x"28",x"1D",x"07",x"4F", -- 0x0AB0
		x"06",x"00",x"21",x"F1",x"0A",x"09",x"7E",x"23", -- 0x0AB8
		x"6E",x"32",x"4C",x"EC",x"7D",x"32",x"4B",x"EC", -- 0x0AC0
		x"3E",x"08",x"32",x"4D",x"EC",x"21",x"14",x"E1", -- 0x0AC8
		x"CB",x"DE",x"C9",x"3A",x"0C",x"E0",x"0F",x"0F", -- 0x0AD0
		x"E6",x"7C",x"C6",x"30",x"6F",x"CD",x"E5",x"0A", -- 0x0AD8
		x"3E",x"E1",x"C3",x"C1",x"0A",x"16",x"02",x"FE", -- 0x0AE0
		x"62",x"D8",x"15",x"FE",x"81",x"D0",x"16",x"03", -- 0x0AE8
		x"C9",x"E1",x"20",x"E1",x"70",x"E1",x"20",x"E1", -- 0x0AF0
		x"70",x"E1",x"20",x"E1",x"02",x"E1",x"34",x"E1", -- 0x0AF8
		x"C0",x"CD",x"8D",x"0C",x"D8",x"16",x"03",x"CD", -- 0x0B00
		x"51",x"0C",x"DA",x"25",x"0B",x"CD",x"A8",x"0C", -- 0x0B08
		x"AF",x"FD",x"77",x"02",x"FD",x"77",x"08",x"FD", -- 0x0B10
		x"77",x"03",x"FD",x"77",x"01",x"32",x"07",x"E1", -- 0x0B18
		x"FD",x"36",x"00",x"C1",x"C9",x"FD",x"36",x"00", -- 0x0B20
		x"00",x"C9",x"3A",x"00",x"EC",x"CB",x"77",x"20", -- 0x0B28
		x"1F",x"CD",x"8D",x"0C",x"D8",x"FD",x"22",x"20", -- 0x0B30
		x"EC",x"3E",x"80",x"FD",x"77",x"0B",x"32",x"11", -- 0x0B38
		x"EC",x"32",x"16",x"EC",x"32",x"1B",x"EC",x"AF", -- 0x0B40
		x"32",x"01",x"EC",x"21",x"00",x"EC",x"CB",x"F6", -- 0x0B48
		x"DD",x"2A",x"20",x"EC",x"3A",x"00",x"EC",x"CB", -- 0x0B50
		x"6F",x"20",x"36",x"DD",x"CB",x"0B",x"7E",x"28", -- 0x0B58
		x"1E",x"DD",x"E5",x"E1",x"01",x"0B",x"00",x"09", -- 0x0B60
		x"E5",x"CD",x"7D",x"0C",x"D1",x"D8",x"7D",x"E6", -- 0x0B68
		x"1F",x"07",x"07",x"12",x"3A",x"01",x"EC",x"3C", -- 0x0B70
		x"32",x"01",x"EC",x"FE",x"04",x"30",x"0D",x"21", -- 0x0B78
		x"11",x"EC",x"CB",x"7E",x"20",x"E2",x"11",x"05", -- 0x0B80
		x"00",x"19",x"18",x"F6",x"21",x"00",x"EC",x"CB", -- 0x0B88
		x"EE",x"DD",x"36",x"01",x"00",x"3A",x"00",x"EC", -- 0x0B90
		x"E6",x"03",x"DD",x"77",x"1D",x"DD",x"77",x"1A", -- 0x0B98
		x"07",x"DD",x"77",x"0D",x"32",x"13",x"EC",x"32", -- 0x0BA0
		x"18",x"EC",x"32",x"1D",x"EC",x"AF",x"DD",x"77", -- 0x0BA8
		x"03",x"DD",x"36",x"00",x"41",x"32",x"01",x"EC", -- 0x0BB0
		x"32",x"00",x"EC",x"C9",x"3A",x"B0",x"E7",x"CB", -- 0x0BB8
		x"77",x"20",x"2A",x"CB",x"67",x"20",x"10",x"AF", -- 0x0BC0
		x"32",x"26",x"E1",x"32",x"36",x"E1",x"3C",x"32", -- 0x0BC8
		x"A9",x"E0",x"21",x"B0",x"E7",x"CB",x"E6",x"CD", -- 0x0BD0
		x"8D",x"0C",x"D8",x"FD",x"22",x"B2",x"E7",x"3E", -- 0x0BD8
		x"80",x"FD",x"77",x"0B",x"AF",x"32",x"B1",x"E7", -- 0x0BE0
		x"21",x"B0",x"E7",x"CB",x"F6",x"DD",x"2A",x"B2", -- 0x0BE8
		x"E7",x"3A",x"B0",x"E7",x"CB",x"6F",x"20",x"28", -- 0x0BF0
		x"3A",x"26",x"E1",x"B7",x"C8",x"3A",x"36",x"E1", -- 0x0BF8
		x"B7",x"C8",x"21",x"90",x"E2",x"11",x"10",x"00", -- 0x0C00
		x"06",x"06",x"7E",x"B7",x"00",x"19",x"10",x"FA", -- 0x0C08
		x"21",x"B0",x"EB",x"06",x"10",x"CB",x"7E",x"C0", -- 0x0C10
		x"23",x"10",x"FA",x"21",x"B0",x"E7",x"CB",x"EE", -- 0x0C18
		x"21",x"B0",x"EB",x"01",x"80",x"10",x"71",x"23", -- 0x0C20
		x"10",x"FC",x"3A",x"B0",x"E7",x"E6",x"03",x"DD", -- 0x0C28
		x"77",x"1D",x"DD",x"77",x"1A",x"07",x"DD",x"77", -- 0x0C30
		x"0D",x"3A",x"B0",x"E7",x"E6",x"08",x"0F",x"0F", -- 0x0C38
		x"F6",x"40",x"DD",x"77",x"01",x"AF",x"DD",x"77", -- 0x0C40
		x"03",x"DD",x"36",x"00",x"41",x"32",x"B0",x"E7", -- 0x0C48
		x"C9",x"21",x"B8",x"EB",x"06",x"02",x"CB",x"4A", -- 0x0C50
		x"28",x"0C",x"21",x"B0",x"EB",x"CB",x"42",x"28", -- 0x0C58
		x"05",x"21",x"A4",x"EB",x"06",x"0C",x"F3",x"CB", -- 0x0C60
		x"7E",x"28",x"0D",x"FB",x"23",x"10",x"F7",x"7A", -- 0x0C68
		x"16",x"03",x"FE",x"03",x"20",x"EB",x"37",x"C9", -- 0x0C70
		x"CB",x"FE",x"FB",x"B7",x"C9",x"21",x"AF",x"EB", -- 0x0C78
		x"06",x"0C",x"F3",x"CB",x"7E",x"28",x"F1",x"FB", -- 0x0C80
		x"2B",x"10",x"F7",x"37",x"C9",x"FD",x"21",x"00", -- 0x0C88
		x"E4",x"06",x"10",x"11",x"30",x"00",x"FD",x"7E", -- 0x0C90
		x"00",x"E6",x"21",x"28",x"06",x"FD",x"19",x"10", -- 0x0C98
		x"F5",x"37",x"C9",x"FD",x"CB",x"00",x"EE",x"C9", -- 0x0CA0
		x"7D",x"07",x"07",x"E6",x"7C",x"FD",x"77",x"0B", -- 0x0CA8
		x"C9",x"3A",x"DF",x"EB",x"0F",x"D2",x"61",x"0E", -- 0x0CB0
		x"E6",x"40",x"C2",x"61",x"0E",x"11",x"E0",x"EB", -- 0x0CB8
		x"2A",x"C4",x"EB",x"CD",x"93",x"0E",x"2A",x"C2", -- 0x0CC0
		x"EB",x"0E",x"20",x"09",x"CB",x"94",x"22",x"C2", -- 0x0CC8
		x"EB",x"2A",x"C4",x"EB",x"7D",x"C6",x"08",x"6F", -- 0x0CD0
		x"22",x"C4",x"EB",x"EB",x"3A",x"A8",x"E0",x"3C", -- 0x0CD8
		x"E6",x"0F",x"32",x"A8",x"E0",x"20",x"28",x"21", -- 0x0CE0
		x"02",x"E1",x"34",x"7E",x"FE",x"10",x"20",x"03", -- 0x0CE8
		x"3E",x"0E",x"77",x"FE",x"02",x"20",x"05",x"3A", -- 0x0CF0
		x"AF",x"E0",x"18",x"0D",x"FE",x"0D",x"20",x"03", -- 0x0CF8
		x"AF",x"18",x"06",x"FE",x"43",x"20",x"08",x"3E", -- 0x0D00
		x"02",x"32",x"D5",x"E0",x"32",x"05",x"C8",x"3E", -- 0x0D08
		x"02",x"2A",x"C0",x"EB",x"F3",x"32",x"06",x"C8", -- 0x0D10
		x"46",x"23",x"4E",x"AF",x"32",x"06",x"C8",x"FB", -- 0x0D18
		x"2B",x"78",x"FE",x"FF",x"20",x"32",x"B9",x"20", -- 0x0D20
		x"2F",x"F3",x"3A",x"D0",x"EB",x"4F",x"2F",x"E6", -- 0x0D28
		x"C0",x"20",x"06",x"79",x"E6",x"BF",x"32",x"D0", -- 0x0D30
		x"EB",x"FB",x"3A",x"02",x"E1",x"FE",x"08",x"30", -- 0x0D38
		x"29",x"21",x"DC",x"98",x"3A",x"02",x"E1",x"B7", -- 0x0D40
		x"CA",x"49",x"0E",x"2A",x"CE",x"EB",x"3D",x"CA", -- 0x0D48
		x"49",x"0E",x"2A",x"C8",x"EB",x"C3",x"49",x"0E", -- 0x0D50
		x"3A",x"D0",x"EB",x"CB",x"77",x"20",x"0B",x"3A", -- 0x0D58
		x"02",x"E1",x"FE",x"44",x"C2",x"49",x"0E",x"C3", -- 0x0D60
		x"67",x"0E",x"3A",x"02",x"E1",x"4F",x"3A",x"D0", -- 0x0D68
		x"EB",x"47",x"E6",x"0F",x"C2",x"C7",x"0D",x"78", -- 0x0D70
		x"CB",x"7F",x"28",x"4B",x"CB",x"77",x"20",x"2C", -- 0x0D78
		x"CB",x"6F",x"20",x"14",x"21",x"D0",x"EB",x"CB", -- 0x0D80
		x"EE",x"CB",x"F6",x"01",x"DC",x"98",x"2A",x"CA", -- 0x0D88
		x"EB",x"ED",x"43",x"CA",x"EB",x"C3",x"49",x"0E", -- 0x0D90
		x"F3",x"3A",x"D0",x"EB",x"F6",x"40",x"32",x"D0", -- 0x0D98
		x"EB",x"FB",x"CB",x"67",x"20",x"06",x"2A",x"CC", -- 0x0DA0
		x"EB",x"C3",x"49",x"0E",x"CB",x"67",x"CA",x"49", -- 0x0DA8
		x"0E",x"3A",x"A8",x"E0",x"FE",x"08",x"C2",x"49", -- 0x0DB0
		x"0E",x"3E",x"42",x"32",x"02",x"E1",x"21",x"D0", -- 0x0DB8
		x"EB",x"CB",x"C6",x"CB",x"CE",x"18",x"48",x"79", -- 0x0DC0
		x"FE",x"43",x"CA",x"19",x"0E",x"CB",x"50",x"20", -- 0x0DC8
		x"78",x"FE",x"42",x"28",x"32",x"CB",x"48",x"C2", -- 0x0DD0
		x"49",x"0E",x"FE",x"41",x"28",x"11",x"CB",x"40", -- 0x0DD8
		x"C2",x"49",x"0E",x"2A",x"CA",x"EB",x"3E",x"40", -- 0x0DE0
		x"32",x"02",x"E1",x"06",x"01",x"18",x"0D",x"3A", -- 0x0DE8
		x"A8",x"E0",x"FE",x"08",x"C2",x"49",x"0E",x"21", -- 0x0DF0
		x"DC",x"98",x"06",x"02",x"F3",x"3A",x"D0",x"EB", -- 0x0DF8
		x"B0",x"32",x"D0",x"EB",x"FB",x"18",x"42",x"3A", -- 0x0E00
		x"A8",x"E0",x"FE",x"08",x"C2",x"49",x"0E",x"21", -- 0x0E08
		x"D0",x"EB",x"CB",x"D6",x"21",x"30",x"80",x"18", -- 0x0E10
		x"30",x"3A",x"A8",x"E0",x"FE",x"08",x"C2",x"49", -- 0x0E18
		x"0E",x"3A",x"99",x"E0",x"B7",x"20",x"22",x"3C", -- 0x0E20
		x"32",x"99",x"E0",x"3E",x"21",x"32",x"9A",x"E0", -- 0x0E28
		x"21",x"E0",x"01",x"22",x"74",x"E1",x"3E",x"01", -- 0x0E30
		x"32",x"76",x"E1",x"32",x"C7",x"E0",x"21",x"D0", -- 0x0E38
		x"EB",x"CB",x"DE",x"21",x"B2",x"80",x"C3",x"49", -- 0x0E40
		x"0E",x"3E",x"02",x"01",x"08",x"00",x"F3",x"32", -- 0x0E48
		x"06",x"C8",x"ED",x"B0",x"AF",x"32",x"06",x"C8", -- 0x0E50
		x"FB",x"22",x"C0",x"EB",x"21",x"DF",x"EB",x"CB", -- 0x0E58
		x"86",x"06",x"02",x"DF",x"C3",x"B1",x"0C",x"AF", -- 0x0E60
		x"32",x"C7",x"EB",x"32",x"02",x"E1",x"3A",x"05", -- 0x0E68
		x"E1",x"3C",x"FE",x"63",x"38",x"02",x"3E",x"63", -- 0x0E70
		x"32",x"05",x"E1",x"21",x"03",x"E1",x"7E",x"3C", -- 0x0E78
		x"FE",x"30",x"38",x"02",x"3E",x"20",x"77",x"32", -- 0x0E80
		x"06",x"E1",x"CD",x"6B",x"19",x"21",x"A6",x"E9", -- 0x0E88
		x"CB",x"FE",x"F7",x"D9",x"21",x"06",x"C8",x"D9", -- 0x0E90
		x"06",x"04",x"C5",x"7E",x"23",x"4E",x"E5",x"6F", -- 0x0E98
		x"79",x"E6",x"0F",x"67",x"79",x"29",x"29",x"29", -- 0x0EA0
		x"01",x"5E",x"99",x"09",x"4F",x"D5",x"CB",x"79", -- 0x0EA8
		x"28",x"03",x"13",x"13",x"13",x"06",x"04",x"D9", -- 0x0EB0
		x"F3",x"36",x"02",x"D9",x"7E",x"12",x"23",x"7E", -- 0x0EB8
		x"D9",x"36",x"00",x"FB",x"D9",x"CB",x"E3",x"CB", -- 0x0EC0
		x"71",x"28",x"02",x"EE",x"20",x"CB",x"79",x"28", -- 0x0EC8
		x"06",x"EE",x"40",x"12",x"1B",x"18",x"02",x"12", -- 0x0ED0
		x"13",x"CB",x"A3",x"23",x"10",x"D9",x"D1",x"21", -- 0x0ED8
		x"04",x"00",x"19",x"EB",x"E1",x"C1",x"23",x"10", -- 0x0EE0
		x"B1",x"C9",x"0E",x"05",x"3A",x"BF",x"EF",x"5F", -- 0x0EE8
		x"04",x"DF",x"06",x"10",x"21",x"E0",x"E0",x"CD", -- 0x0EF0
		x"13",x"0F",x"10",x"FB",x"D9",x"11",x"01",x"00", -- 0x0EF8
		x"2A",x"0C",x"E0",x"19",x"22",x"0C",x"E0",x"1D", -- 0x0F00
		x"2A",x"0E",x"E0",x"ED",x"5A",x"22",x"0E",x"E0", -- 0x0F08
		x"D9",x"18",x"DD",x"79",x"B7",x"28",x"04",x"34", -- 0x0F10
		x"2C",x"0D",x"C9",x"7B",x"B7",x"20",x"03",x"35", -- 0x0F18
		x"18",x"11",x"3D",x"20",x"04",x"CB",x"06",x"18", -- 0x0F20
		x"0A",x"3D",x"20",x"04",x"CB",x"0E",x"18",x"03", -- 0x0F28
		x"7E",x"2F",x"77",x"2C",x"3A",x"0C",x"E0",x"E6", -- 0x0F30
		x"0F",x"3C",x"4F",x"0F",x"E6",x"03",x"5F",x"C9", -- 0x0F38
		x"21",x"20",x"E0",x"AF",x"BE",x"28",x"0E",x"1E", -- 0x0F40
		x"01",x"E5",x"CD",x"5A",x"0F",x"06",x"04",x"DF", -- 0x0F48
		x"CD",x"62",x"0F",x"E1",x"35",x"06",x"04",x"DF", -- 0x0F50
		x"18",x"E6",x"7B",x"21",x"D4",x"E0",x"F3",x"B6", -- 0x0F58
		x"18",x"07",x"21",x"D4",x"E0",x"7B",x"2F",x"F3", -- 0x0F60
		x"A6",x"77",x"32",x"04",x"C8",x"FB",x"C9",x"AF", -- 0x0F68
		x"32",x"28",x"E0",x"CD",x"8D",x"11",x"3E",x"80", -- 0x0F70
		x"32",x"01",x"E0",x"0E",x"0F",x"CD",x"78",x"11", -- 0x0F78
		x"0E",x"00",x"CD",x"78",x"11",x"0E",x"10",x"CD", -- 0x0F80
		x"78",x"11",x"AF",x"32",x"00",x"E0",x"32",x"01", -- 0x0F88
		x"E0",x"CD",x"E7",x"2C",x"CD",x"FD",x"2C",x"CD", -- 0x0F90
		x"A7",x"02",x"CD",x"B6",x"11",x"CD",x"E0",x"11", -- 0x0F98
		x"CD",x"89",x"18",x"21",x"28",x"E0",x"34",x"7E", -- 0x0FA0
		x"0F",x"D2",x"75",x"10",x"DD",x"21",x"B7",x"A1", -- 0x0FA8
		x"CD",x"CC",x"2C",x"CD",x"9C",x"12",x"CD",x"F3", -- 0x0FB0
		x"11",x"CD",x"6C",x"11",x"CD",x"22",x"11",x"21", -- 0x0FB8
		x"00",x"72",x"22",x"2B",x"E0",x"2A",x"00",x"72", -- 0x0FC0
		x"22",x"29",x"E0",x"AF",x"6F",x"67",x"22",x"02", -- 0x0FC8
		x"E1",x"32",x"06",x"E1",x"3A",x"02",x"E0",x"E6", -- 0x0FD0
		x"02",x"CA",x"06",x"10",x"0E",x"03",x"C5",x"21", -- 0x0FD8
		x"0A",x"11",x"11",x"5C",x"EB",x"01",x"08",x"00", -- 0x0FE0
		x"ED",x"B0",x"C1",x"06",x"20",x"CD",x"55",x"10", -- 0x0FE8
		x"06",x"28",x"DF",x"0D",x"79",x"B7",x"28",x"54", -- 0x0FF0
		x"21",x"00",x"00",x"22",x"5D",x"EB",x"22",x"61", -- 0x0FF8
		x"EB",x"06",x"08",x"DF",x"18",x"D8",x"21",x"12", -- 0x1000
		x"11",x"11",x"5C",x"EB",x"01",x"08",x"00",x"ED", -- 0x1008
		x"B0",x"06",x"38",x"CD",x"55",x"10",x"06",x"18", -- 0x1010
		x"CD",x"65",x"10",x"21",x"00",x"00",x"22",x"5D", -- 0x1018
		x"EB",x"22",x"61",x"EB",x"21",x"1A",x"11",x"11", -- 0x1020
		x"00",x"EB",x"01",x"04",x"00",x"ED",x"B0",x"06", -- 0x1028
		x"30",x"DF",x"01",x"FF",x"04",x"C5",x"06",x"01", -- 0x1030
		x"DF",x"C1",x"79",x"3C",x"E6",x"03",x"4F",x"5F", -- 0x1038
		x"16",x"00",x"21",x"1E",x"11",x"19",x"7E",x"32", -- 0x1040
		x"00",x"EB",x"10",x"E9",x"06",x"A0",x"DF",x"06", -- 0x1048
		x"00",x"DF",x"C3",x"AA",x"10",x"C5",x"21",x"5E", -- 0x1050
		x"EB",x"35",x"21",x"62",x"EB",x"34",x"06",x"02", -- 0x1058
		x"DF",x"C1",x"10",x"F1",x"C9",x"C5",x"21",x"5E", -- 0x1060
		x"EB",x"34",x"21",x"62",x"EB",x"35",x"06",x"02", -- 0x1068
		x"DF",x"C1",x"10",x"F1",x"C9",x"DD",x"21",x"16", -- 0x1070
		x"A3",x"CD",x"CC",x"2C",x"CD",x"9C",x"12",x"21", -- 0x1078
		x"92",x"D0",x"CD",x"6F",x"11",x"21",x"EA",x"A4", -- 0x1080
		x"CD",x"22",x"02",x"CD",x"46",x"6C",x"21",x"5D", -- 0x1088
		x"73",x"22",x"2B",x"E0",x"2A",x"5D",x"73",x"22", -- 0x1090
		x"29",x"E0",x"21",x"03",x"01",x"22",x"02",x"E1", -- 0x1098
		x"7C",x"32",x"06",x"E1",x"06",x"00",x"DF",x"06", -- 0x10A0
		x"78",x"DF",x"CD",x"A7",x"02",x"CD",x"B6",x"11", -- 0x10A8
		x"CD",x"9C",x"12",x"DD",x"21",x"00",x"E1",x"CD", -- 0x10B0
		x"23",x"19",x"CD",x"22",x"12",x"2A",x"02",x"E0", -- 0x10B8
		x"23",x"22",x"02",x"E0",x"DD",x"21",x"FF",x"A1", -- 0x10C0
		x"CD",x"CC",x"2C",x"21",x"28",x"E0",x"7E",x"0F", -- 0x10C8
		x"D4",x"22",x"11",x"3E",x"0C",x"EF",x"21",x"E0", -- 0x10D0
		x"E0",x"06",x"10",x"CD",x"13",x"2D",x"21",x"FF", -- 0x10D8
		x"FF",x"22",x"04",x"E1",x"AF",x"6F",x"67",x"22", -- 0x10E0
		x"0C",x"E0",x"22",x"0E",x"E0",x"32",x"2D",x"E0", -- 0x10E8
		x"32",x"45",x"EC",x"32",x"19",x"E1",x"3C",x"32", -- 0x10F0
		x"A6",x"E0",x"3C",x"32",x"00",x"E1",x"06",x"01", -- 0x10F8
		x"DF",x"3E",x"0C",x"01",x"EA",x"0E",x"FF",x"C3", -- 0x1100
		x"FB",x"14",x"D0",x"46",x"81",x"20",x"D2",x"46", -- 0x1108
		x"61",x"20",x"6C",x"A6",x"81",x"20",x"6C",x"A6", -- 0x1110
		x"41",x"20",x"6C",x"A6",x"61",x"20",x"68",x"68", -- 0x1118
		x"64",x"64",x"3E",x"0D",x"01",x"29",x"11",x"FF", -- 0x1120
		x"C9",x"06",x"14",x"DF",x"21",x"96",x"A4",x"CD", -- 0x1128
		x"22",x"02",x"06",x"3C",x"DF",x"3A",x"97",x"A4", -- 0x1130
		x"47",x"2A",x"98",x"A4",x"CD",x"47",x"02",x"18", -- 0x1138
		x"E8",x"3A",x"2A",x"E0",x"4F",x"21",x"29",x"E0", -- 0x1140
		x"35",x"C0",x"2A",x"2B",x"E0",x"7E",x"B7",x"20", -- 0x1148
		x"0D",x"3A",x"28",x"E0",x"0F",x"21",x"00",x"72", -- 0x1150
		x"38",x"03",x"21",x"5D",x"73",x"7E",x"32",x"29", -- 0x1158
		x"E0",x"23",x"7E",x"32",x"2A",x"E0",x"4F",x"23", -- 0x1160
		x"22",x"2B",x"E0",x"C9",x"21",x"90",x"D0",x"11", -- 0x1168
		x"44",x"A3",x"01",x"06",x"17",x"C3",x"75",x"02", -- 0x1170
		x"3A",x"00",x"E0",x"E6",x"80",x"C8",x"F3",x"2A", -- 0x1178
		x"22",x"E2",x"71",x"23",x"7D",x"E6",x"1F",x"6F", -- 0x1180
		x"22",x"22",x"E2",x"FB",x"C9",x"CD",x"A2",x"11", -- 0x1188
		x"AF",x"67",x"6F",x"22",x"D2",x"E0",x"22",x"D5", -- 0x1190
		x"E0",x"22",x"02",x"C8",x"22",x"05",x"C8",x"C3", -- 0x1198
		x"08",x"2D",x"21",x"D4",x"E0",x"3A",x"04",x"C0", -- 0x11A0
		x"E6",x"10",x"28",x"05",x"CB",x"BE",x"C3",x"08", -- 0x11A8
		x"2D",x"CB",x"FE",x"C3",x"08",x"2D",x"21",x"40", -- 0x11B0
		x"D0",x"01",x"80",x"03",x"CD",x"E0",x"01",x"21", -- 0x11B8
		x"40",x"D4",x"01",x"80",x"03",x"16",x"00",x"C3", -- 0x11C0
		x"E2",x"01",x"21",x"40",x"D0",x"01",x"1D",x"1C", -- 0x11C8
		x"16",x"30",x"CD",x"53",x"02",x"21",x"40",x"D4", -- 0x11D0
		x"01",x"1D",x"1C",x"16",x"00",x"C3",x"53",x"02", -- 0x11D8
		x"21",x"01",x"D8",x"16",x"F8",x"CD",x"ED",x"11", -- 0x11E0
		x"21",x"11",x"D8",x"16",x"80",x"01",x"0E",x"20", -- 0x11E8
		x"C3",x"53",x"02",x"21",x"22",x"D5",x"01",x"02", -- 0x11F0
		x"0E",x"3E",x"02",x"21",x"46",x"A4",x"C3",x"22", -- 0x11F8
		x"02",x"3A",x"00",x"E0",x"0F",x"D8",x"21",x"E0", -- 0x1200
		x"A4",x"CD",x"22",x"02",x"3A",x"00",x"E0",x"0F", -- 0x1208
		x"D8",x"0E",x"00",x"C3",x"14",x"13",x"06",x"02", -- 0x1210
		x"11",x"11",x"E0",x"F3",x"CD",x"0E",x"02",x"FB", -- 0x1218
		x"18",x"EA",x"21",x"40",x"D4",x"01",x"31",x"16", -- 0x1220
		x"CD",x"49",x"02",x"21",x"40",x"D0",x"3A",x"01", -- 0x1228
		x"E1",x"B7",x"06",x"16",x"28",x"32",x"11",x"20", -- 0x1230
		x"00",x"0E",x"42",x"D9",x"4F",x"11",x"64",x"00", -- 0x1238
		x"CD",x"86",x"12",x"CD",x"8E",x"12",x"11",x"0A", -- 0x1240
		x"00",x"CD",x"86",x"12",x"CD",x"8E",x"12",x"D9", -- 0x1248
		x"C5",x"D5",x"E5",x"11",x"00",x"04",x"19",x"11", -- 0x1250
		x"20",x"00",x"36",x"32",x"19",x"10",x"FB",x"E1", -- 0x1258
		x"D1",x"C1",x"D9",x"51",x"CD",x"8E",x"12",x"D9", -- 0x1260
		x"0E",x"30",x"C3",x"49",x"02",x"21",x"40",x"D4", -- 0x1268
		x"01",x"31",x"16",x"CD",x"49",x"02",x"21",x"40", -- 0x1270
		x"D0",x"3A",x"01",x"E1",x"06",x"16",x"B7",x"28", -- 0x1278
		x"E7",x"3D",x"28",x"E4",x"18",x"B0",x"79",x"BB", -- 0x1280
		x"D8",x"93",x"4F",x"14",x"18",x"F9",x"7A",x"B7", -- 0x1288
		x"D9",x"28",x"06",x"71",x"19",x"05",x"3D",x"20", -- 0x1290
		x"FA",x"0D",x"D9",x"C9",x"21",x"5E",x"D4",x"01", -- 0x1298
		x"33",x"1C",x"CD",x"49",x"02",x"21",x"5F",x"D4", -- 0x12A0
		x"01",x"19",x"1C",x"CD",x"49",x"02",x"21",x"7F", -- 0x12A8
		x"D5",x"01",x"1A",x"0A",x"CD",x"49",x"02",x"21", -- 0x12B0
		x"C6",x"A4",x"CD",x"22",x"02",x"0E",x"05",x"CD", -- 0x12B8
		x"14",x"13",x"0E",x"0A",x"CD",x"14",x"13",x"3A", -- 0x12C0
		x"01",x"E0",x"07",x"D0",x"0E",x"0F",x"C3",x"14", -- 0x12C8
		x"13",x"3A",x"00",x"E0",x"07",x"D0",x"3A",x"00", -- 0x12D0
		x"E1",x"E6",x"01",x"11",x"57",x"E0",x"3E",x"0F", -- 0x12D8
		x"20",x"05",x"11",x"4F",x"E0",x"3E",x"0A",x"F5", -- 0x12E0
		x"06",x"08",x"CD",x"FA",x"01",x"F1",x"4F",x"CD", -- 0x12E8
		x"14",x"13",x"3A",x"00",x"E1",x"E6",x"01",x"11", -- 0x12F0
		x"50",x"E0",x"20",x"03",x"11",x"48",x"E0",x"06", -- 0x12F8
		x"08",x"21",x"40",x"E0",x"D5",x"CD",x"77",x"6B", -- 0x1300
		x"E1",x"D8",x"11",x"40",x"E0",x"01",x"08",x"00", -- 0x1308
		x"ED",x"B0",x"0E",x"05",x"06",x"00",x"21",x"32", -- 0x1310
		x"13",x"09",x"5E",x"23",x"56",x"23",x"D5",x"5E", -- 0x1318
		x"23",x"56",x"23",x"46",x"E1",x"78",x"07",x"D2", -- 0x1320
		x"EE",x"01",x"06",x"07",x"CD",x"63",x"02",x"AF", -- 0x1328
		x"77",x"C9",x"80",x"D3",x"10",x"E0",x"02",x"9E", -- 0x1330
		x"D1",x"40",x"E0",x"88",x"5E",x"D0",x"48",x"E0", -- 0x1338
		x"88",x"BE",x"D2",x"50",x"E0",x"88",x"3E",x"80", -- 0x1340
		x"32",x"00",x"E0",x"AF",x"32",x"C7",x"EB",x"3E", -- 0x1348
		x"0C",x"01",x"EA",x"0E",x"FF",x"CD",x"A2",x"11", -- 0x1350
		x"CD",x"08",x"2D",x"CD",x"A7",x"02",x"CD",x"E0", -- 0x1358
		x"11",x"CD",x"E7",x"2C",x"CD",x"B6",x"11",x"2A", -- 0x1360
		x"10",x"E0",x"7D",x"B4",x"3A",x"00",x"E0",x"C2", -- 0x1368
		x"77",x"13",x"E6",x"04",x"CA",x"6F",x"0F",x"DD", -- 0x1370
		x"21",x"E0",x"A1",x"E6",x"04",x"28",x"04",x"DD", -- 0x1378
		x"21",x"BA",x"A2",x"CD",x"B6",x"11",x"CD",x"CC", -- 0x1380
		x"2C",x"DD",x"21",x"00",x"E1",x"CD",x"23",x"19", -- 0x1388
		x"CD",x"9C",x"12",x"CD",x"22",x"12",x"CD",x"01", -- 0x1390
		x"12",x"3A",x"00",x"E0",x"E6",x"04",x"20",x"0B", -- 0x1398
		x"CD",x"6C",x"11",x"21",x"46",x"A4",x"CD",x"22", -- 0x13A0
		x"02",x"18",x"1C",x"21",x"52",x"A5",x"CD",x"22", -- 0x13A8
		x"02",x"21",x"01",x"00",x"22",x"98",x"E0",x"3E", -- 0x13B0
		x"1E",x"32",x"9A",x"E0",x"CD",x"42",x"17",x"2A", -- 0x13B8
		x"10",x"E0",x"7D",x"B4",x"CC",x"22",x"11",x"06", -- 0x13C0
		x"02",x"DF",x"2A",x"10",x"E0",x"7D",x"B4",x"28", -- 0x13C8
		x"41",x"21",x"58",x"A4",x"3A",x"00",x"E0",x"E6", -- 0x13D0
		x"04",x"28",x"16",x"3A",x"F4",x"EF",x"B7",x"28", -- 0x13D8
		x"13",x"3E",x"0D",x"EF",x"21",x"4A",x"D1",x"01", -- 0x13E0
		x"01",x"0B",x"16",x"30",x"CD",x"53",x"02",x"18", -- 0x13E8
		x"03",x"CD",x"22",x"02",x"2A",x"10",x"E0",x"7D", -- 0x13F0
		x"6C",x"67",x"11",x"FE",x"FF",x"19",x"38",x"61", -- 0x13F8
		x"21",x"6D",x"A4",x"3A",x"00",x"E0",x"E6",x"04", -- 0x1400
		x"CC",x"22",x"02",x"3A",x"00",x"C0",x"E6",x"01", -- 0x1408
		x"28",x"45",x"3A",x"00",x"E0",x"E6",x"04",x"CA", -- 0x1410
		x"C7",x"13",x"2A",x"98",x"E0",x"7D",x"B4",x"20", -- 0x1418
		x"1C",x"21",x"9A",x"E0",x"35",x"C2",x"C7",x"13", -- 0x1420
		x"21",x"00",x"E0",x"CB",x"96",x"3E",x"0D",x"EF", -- 0x1428
		x"2A",x"98",x"A4",x"3A",x"97",x"A4",x"47",x"CD", -- 0x1430
		x"47",x"02",x"C3",x"67",x"13",x"21",x"9A",x"E0", -- 0x1438
		x"35",x"C2",x"C7",x"13",x"36",x"1E",x"21",x"C4", -- 0x1440
		x"78",x"11",x"99",x"E0",x"06",x"02",x"CD",x"0E", -- 0x1448
		x"02",x"CD",x"42",x"17",x"C3",x"C7",x"13",x"21", -- 0x1450
		x"C4",x"78",x"CD",x"16",x"12",x"3E",x"01",x"18", -- 0x1458
		x"1A",x"21",x"80",x"A4",x"3A",x"00",x"E0",x"E6", -- 0x1460
		x"04",x"CC",x"22",x"02",x"3A",x"00",x"C0",x"E6", -- 0x1468
		x"02",x"20",x"98",x"21",x"C6",x"78",x"CD",x"16", -- 0x1470
		x"12",x"3E",x"83",x"32",x"01",x"E0",x"3E",x"0D", -- 0x1478
		x"EF",x"2A",x"98",x"A4",x"3A",x"97",x"A4",x"47", -- 0x1480
		x"CD",x"47",x"02",x"3A",x"01",x"C0",x"2F",x"E6", -- 0x1488
		x"30",x"B7",x"C4",x"67",x"17",x"4F",x"3A",x"00", -- 0x1490
		x"E1",x"B1",x"32",x"00",x"E1",x"3A",x"02",x"C0", -- 0x1498
		x"2F",x"E6",x"30",x"C4",x"67",x"17",x"4F",x"3A", -- 0x14A0
		x"80",x"E1",x"B1",x"32",x"80",x"E1",x"21",x"48", -- 0x14A8
		x"E0",x"01",x"30",x"00",x"50",x"CD",x"E2",x"01", -- 0x14B0
		x"3A",x"00",x"E0",x"E6",x"04",x"F6",x"80",x"32", -- 0x14B8
		x"00",x"E0",x"2A",x"04",x"E0",x"23",x"22",x"04", -- 0x14C0
		x"E0",x"CD",x"9C",x"12",x"2A",x"03",x"C0",x"7D", -- 0x14C8
		x"E6",x"07",x"28",x"05",x"7C",x"E6",x"07",x"20", -- 0x14D0
		x"06",x"21",x"00",x"02",x"22",x"10",x"E0",x"CD", -- 0x14D8
		x"A2",x"11",x"CD",x"89",x"18",x"CD",x"91",x"18", -- 0x14E0
		x"3E",x"01",x"32",x"A6",x"E0",x"3E",x"83",x"32", -- 0x14E8
		x"00",x"E0",x"CD",x"A7",x"02",x"CD",x"B6",x"11", -- 0x14F0
		x"CD",x"08",x"2D",x"CD",x"90",x"11",x"AF",x"32", -- 0x14F8
		x"C7",x"EB",x"0E",x"00",x"CD",x"78",x"11",x"0E", -- 0x1500
		x"10",x"CD",x"78",x"11",x"21",x"00",x"E4",x"01", -- 0x1508
		x"00",x"03",x"16",x"00",x"CD",x"E2",x"01",x"AF", -- 0x1510
		x"32",x"A8",x"E0",x"3A",x"02",x"E1",x"FE",x"09", -- 0x1518
		x"38",x"02",x"3E",x"09",x"32",x"02",x"E1",x"3E", -- 0x1520
		x"01",x"F3",x"32",x"06",x"C8",x"3A",x"06",x"E1", -- 0x1528
		x"32",x"03",x"E1",x"E6",x"3F",x"21",x"00",x"80", -- 0x1530
		x"CD",x"36",x"19",x"3A",x"02",x"E1",x"B7",x"28", -- 0x1538
		x"11",x"47",x"7E",x"FE",x"FD",x"28",x"08",x"CB", -- 0x1540
		x"7E",x"20",x"01",x"23",x"23",x"18",x"F3",x"23", -- 0x1548
		x"10",x"F0",x"22",x"A0",x"E9",x"AF",x"32",x"06", -- 0x1550
		x"C8",x"FB",x"AF",x"6F",x"67",x"22",x"78",x"E0", -- 0x1558
		x"22",x"7A",x"E0",x"22",x"7C",x"E0",x"22",x"7E", -- 0x1560
		x"E0",x"22",x"90",x"E0",x"32",x"92",x"E0",x"32", -- 0x1568
		x"93",x"E0",x"22",x"94",x"E0",x"32",x"96",x"E0", -- 0x1570
		x"22",x"14",x"E1",x"22",x"7C",x"E1",x"22",x"7E", -- 0x1578
		x"E1",x"32",x"A1",x"E0",x"32",x"18",x"E1",x"22", -- 0x1580
		x"B0",x"E7",x"32",x"A2",x"E0",x"32",x"07",x"E1", -- 0x1588
		x"32",x"17",x"E1",x"32",x"C2",x"E0",x"32",x"B4", -- 0x1590
		x"E7",x"32",x"1E",x"E1",x"32",x"49",x"EC",x"32", -- 0x1598
		x"48",x"EC",x"32",x"1D",x"E1",x"32",x"1B",x"E1", -- 0x15A0
		x"32",x"EA",x"E7",x"32",x"A5",x"E0",x"32",x"6B", -- 0x15A8
		x"E1",x"32",x"70",x"E1",x"32",x"16",x"E1",x"32", -- 0x15B0
		x"F0",x"E3",x"32",x"A4",x"E0",x"32",x"C7",x"E0", -- 0x15B8
		x"32",x"91",x"E7",x"32",x"1A",x"E1",x"32",x"A9", -- 0x15C0
		x"E0",x"3C",x"32",x"C5",x"E0",x"3C",x"32",x"AD", -- 0x15C8
		x"E0",x"3A",x"1F",x"E1",x"E6",x"03",x"32",x"1F", -- 0x15D0
		x"E1",x"3E",x"28",x"32",x"AE",x"E0",x"3A",x"03", -- 0x15D8
		x"E1",x"FE",x"20",x"3E",x"03",x"38",x"02",x"3E", -- 0x15E0
		x"04",x"32",x"9B",x"E0",x"CD",x"40",x"19",x"21", -- 0x15E8
		x"00",x"E3",x"06",x"0F",x"11",x"10",x"00",x"CD", -- 0x15F0
		x"48",x"19",x"3A",x"07",x"EC",x"F5",x"21",x"00", -- 0x15F8
		x"EC",x"01",x"60",x"00",x"50",x"CD",x"E2",x"01", -- 0x1600
		x"F1",x"32",x"07",x"EC",x"3E",x"80",x"32",x"11", -- 0x1608
		x"EC",x"32",x"16",x"EC",x"32",x"1B",x"EC",x"21", -- 0x1610
		x"A0",x"EB",x"01",x"20",x"00",x"50",x"CD",x"E2", -- 0x1618
		x"01",x"DD",x"21",x"20",x"E1",x"CD",x"49",x"18", -- 0x1620
		x"DD",x"21",x"30",x"E1",x"CD",x"49",x"18",x"21", -- 0x1628
		x"E0",x"E7",x"01",x"1F",x"00",x"16",x"00",x"CD", -- 0x1630
		x"E2",x"01",x"21",x"F0",x"E7",x"22",x"E8",x"E7", -- 0x1638
		x"3E",x"0A",x"32",x"ED",x"E7",x"CD",x"4D",x"07", -- 0x1640
		x"3E",x"07",x"32",x"4E",x"EC",x"CD",x"3F",x"0A", -- 0x1648
		x"21",x"A0",x"EB",x"16",x"83",x"0E",x"04",x"CD", -- 0x1650
		x"E2",x"01",x"21",x"B4",x"A8",x"22",x"58",x"E1", -- 0x1658
		x"3E",x"70",x"32",x"63",x"E1",x"3E",x"E0",x"32", -- 0x1660
		x"46",x"E1",x"21",x"14",x"A8",x"CD",x"70",x"17", -- 0x1668
		x"3A",x"03",x"E1",x"E6",x"1F",x"4F",x"09",x"7E", -- 0x1670
		x"32",x"78",x"E1",x"3E",x"05",x"32",x"79",x"E1", -- 0x1678
		x"3C",x"32",x"F1",x"E9",x"21",x"9C",x"A8",x"CD", -- 0x1680
		x"70",x"17",x"3A",x"03",x"E1",x"E6",x"18",x"0F", -- 0x1688
		x"0F",x"0F",x"4F",x"06",x"00",x"09",x"7E",x"32", -- 0x1690
		x"F0",x"E9",x"CD",x"44",x"2B",x"CD",x"68",x"2B", -- 0x1698
		x"AF",x"32",x"05",x"EC",x"3A",x"53",x"E1",x"32", -- 0x16A0
		x"54",x"E1",x"CD",x"8A",x"2B",x"3E",x"01",x"32", -- 0x16A8
		x"76",x"E1",x"21",x"F0",x"00",x"22",x"74",x"E1", -- 0x16B0
		x"DD",x"21",x"60",x"E2",x"2E",x"04",x"11",x"10", -- 0x16B8
		x"00",x"01",x"58",x"E0",x"06",x"03",x"DD",x"75", -- 0x16C0
		x"0B",x"7D",x"C6",x"04",x"6F",x"DD",x"71",x"08", -- 0x16C8
		x"79",x"C6",x"08",x"4F",x"DD",x"19",x"10",x"EE", -- 0x16D0
		x"21",x"48",x"68",x"11",x"04",x"04",x"06",x"06", -- 0x16D8
		x"DD",x"75",x"04",x"DD",x"74",x"05",x"19",x"C5", -- 0x16E0
		x"01",x"10",x"00",x"DD",x"09",x"C1",x"10",x"F0", -- 0x16E8
		x"CD",x"9C",x"12",x"CD",x"4E",x"19",x"CD",x"22", -- 0x16F0
		x"12",x"21",x"00",x"D7",x"01",x"05",x"06",x"CD", -- 0x16F8
		x"49",x"02",x"CD",x"67",x"18",x"3A",x"00",x"E1", -- 0x1700
		x"CB",x"6F",x"CC",x"65",x"19",x"3E",x"50",x"32", -- 0x1708
		x"C1",x"E0",x"3A",x"02",x"E1",x"B7",x"20",x"0E", -- 0x1710
		x"6F",x"67",x"22",x"55",x"E1",x"32",x"57",x"E1", -- 0x1718
		x"22",x"65",x"E1",x"32",x"67",x"E1",x"CD",x"6D", -- 0x1720
		x"12",x"DD",x"21",x"E8",x"1A",x"CD",x"19",x"2D", -- 0x1728
		x"3E",x"20",x"32",x"DE",x"EB",x"21",x"DF",x"EB", -- 0x1730
		x"36",x"00",x"21",x"C7",x"EB",x"36",x"01",x"C3", -- 0x1738
		x"F5",x"1A",x"3A",x"98",x"E0",x"DD",x"21",x"B8", -- 0x1740
		x"D1",x"CD",x"53",x"17",x"3A",x"99",x"E0",x"DD", -- 0x1748
		x"21",x"18",x"D2",x"07",x"07",x"C6",x"80",x"DD", -- 0x1750
		x"77",x"00",x"3C",x"DD",x"77",x"01",x"3C",x"DD", -- 0x1758
		x"77",x"20",x"3C",x"DD",x"77",x"21",x"C9",x"3A", -- 0x1760
		x"00",x"E0",x"E6",x"04",x"C8",x"3E",x"10",x"C9", -- 0x1768
		x"3A",x"04",x"C0",x"E6",x"60",x"0F",x"0F",x"0F", -- 0x1770
		x"0F",x"4F",x"06",x"00",x"09",x"7E",x"23",x"66", -- 0x1778
		x"6F",x"C9",x"21",x"41",x"D0",x"01",x"1D",x"1C", -- 0x1780
		x"16",x"30",x"CD",x"53",x"02",x"3E",x"01",x"32", -- 0x1788
		x"C4",x"E0",x"3A",x"00",x"E0",x"07",x"D2",x"20", -- 0x1790
		x"18",x"DD",x"21",x"43",x"A2",x"CD",x"CC",x"2C", -- 0x1798
		x"3A",x"02",x"E1",x"B7",x"CC",x"28",x"18",x"3A", -- 0x17A0
		x"03",x"E1",x"E6",x"1F",x"4F",x"3E",x"20",x"91", -- 0x17A8
		x"FE",x"01",x"21",x"47",x"A6",x"28",x"1F",x"06", -- 0x17B0
		x"00",x"FE",x"0A",x"38",x"05",x"D6",x"0A",x"04", -- 0x17B8
		x"18",x"F7",x"4F",x"C5",x"21",x"55",x"A6",x"CD", -- 0x17C0
		x"22",x"02",x"C1",x"78",x"32",x"D1",x"D1",x"79", -- 0x17C8
		x"32",x"F1",x"D1",x"21",x"5D",x"A6",x"CD",x"22", -- 0x17D0
		x"02",x"21",x"48",x"D4",x"16",x"3C",x"01",x"08", -- 0x17D8
		x"1C",x"CD",x"53",x"02",x"21",x"BD",x"A4",x"CD", -- 0x17E0
		x"22",x"02",x"CD",x"2F",x"2D",x"21",x"B1",x"A4", -- 0x17E8
		x"20",x"03",x"21",x"A5",x"A4",x"CD",x"22",x"02", -- 0x17F0
		x"06",x"DC",x"DF",x"2A",x"A7",x"A4",x"01",x"03", -- 0x17F8
		x"08",x"16",x"30",x"CD",x"53",x"02",x"21",x"50", -- 0x1800
		x"D0",x"01",x"0D",x"1C",x"CD",x"53",x"02",x"0E", -- 0x1808
		x"02",x"C5",x"06",x"33",x"DF",x"C1",x"0D",x"20", -- 0x1810
		x"F8",x"0E",x"11",x"CD",x"78",x"11",x"18",x"03", -- 0x1818
		x"CD",x"F3",x"11",x"AF",x"32",x"C4",x"E0",x"F7", -- 0x1820
		x"3A",x"03",x"E1",x"E6",x"03",x"FE",x"03",x"21", -- 0x1828
		x"2B",x"A6",x"CC",x"22",x"02",x"21",x"17",x"A7", -- 0x1830
		x"3A",x"03",x"E1",x"0F",x"E6",x"0E",x"4F",x"06", -- 0x1838
		x"00",x"09",x"7E",x"23",x"66",x"6F",x"C3",x"22", -- 0x1840
		x"02",x"DD",x"7E",x"00",x"E6",x"E3",x"DD",x"77", -- 0x1848
		x"00",x"E6",x"8E",x"FE",x"82",x"C0",x"DD",x"7E", -- 0x1850
		x"0B",x"E6",x"7C",x"0F",x"0F",x"4F",x"06",x"00", -- 0x1858
		x"21",x"A0",x"EB",x"09",x"36",x"80",x"C9",x"21", -- 0x1860
		x"A0",x"D3",x"11",x"E0",x"FF",x"0E",x"30",x"06", -- 0x1868
		x"06",x"3A",x"9B",x"E0",x"B7",x"28",x"0D",x"0E", -- 0x1870
		x"68",x"71",x"19",x"05",x"3D",x"20",x"FA",x"78", -- 0x1878
		x"B7",x"C8",x"0E",x"30",x"71",x"19",x"10",x"FC", -- 0x1880
		x"C9",x"DD",x"21",x"00",x"E1",x"1E",x"00",x"18", -- 0x1888
		x"06",x"DD",x"21",x"80",x"E1",x"1E",x"01",x"DD", -- 0x1890
		x"7E",x"03",x"FE",x"1F",x"38",x"04",x"DD",x"CB", -- 0x1898
		x"00",x"A6",x"DD",x"E5",x"E1",x"01",x"80",x"00", -- 0x18A0
		x"50",x"DD",x"CB",x"00",x"66",x"CC",x"E2",x"01", -- 0x18A8
		x"21",x"00",x"08",x"3A",x"03",x"C0",x"E6",x"10", -- 0x18B0
		x"20",x"03",x"21",x"01",x"00",x"DD",x"75",x"10", -- 0x18B8
		x"DD",x"74",x"11",x"AF",x"32",x"07",x"EC",x"DD", -- 0x18C0
		x"CB",x"00",x"66",x"20",x"1C",x"DD",x"36",x"0A", -- 0x18C8
		x"02",x"DD",x"77",x"40",x"DD",x"77",x"41",x"DD", -- 0x18D0
		x"77",x"02",x"DD",x"77",x"14",x"DD",x"77",x"15", -- 0x18D8
		x"DD",x"77",x"16",x"DD",x"77",x"13",x"DD",x"77", -- 0x18E0
		x"6A",x"DD",x"77",x"19",x"DD",x"77",x"1F",x"DD", -- 0x18E8
		x"77",x"64",x"DD",x"77",x"5D",x"DD",x"77",x"5E", -- 0x18F0
		x"DD",x"77",x"5F",x"DD",x"77",x"4D",x"DD",x"77", -- 0x18F8
		x"4E",x"DD",x"77",x"4F",x"DD",x"77",x"55",x"DD", -- 0x1900
		x"77",x"56",x"DD",x"77",x"57",x"DD",x"77",x"65", -- 0x1908
		x"DD",x"77",x"66",x"DD",x"77",x"67",x"DD",x"77", -- 0x1910
		x"20",x"DD",x"77",x"30",x"DD",x"36",x"04",x"C8", -- 0x1918
		x"DD",x"73",x"00",x"21",x"80",x"78",x"3A",x"03", -- 0x1920
		x"C0",x"07",x"07",x"E6",x"03",x"4F",x"06",x"00", -- 0x1928
		x"09",x"7E",x"DD",x"77",x"01",x"C9",x"07",x"4F", -- 0x1930
		x"06",x"00",x"09",x"7E",x"23",x"66",x"6F",x"C9", -- 0x1938
		x"21",x"60",x"E2",x"06",x"09",x"11",x"10",x"00", -- 0x1940
		x"AF",x"77",x"19",x"10",x"FC",x"C9",x"3A",x"00", -- 0x1948
		x"E0",x"07",x"D0",x"3A",x"00",x"E1",x"21",x"9F", -- 0x1950
		x"D4",x"0F",x"38",x"03",x"21",x"3F",x"D7",x"01", -- 0x1958
		x"00",x"03",x"C3",x"49",x"02",x"CD",x"E0",x"11", -- 0x1960
		x"3A",x"03",x"E1",x"F5",x"3C",x"E6",x"07",x"FE", -- 0x1968
		x"07",x"3E",x"00",x"20",x"08",x"21",x"5C",x"98", -- 0x1970
		x"22",x"CC",x"EB",x"3E",x"80",x"32",x"D0",x"EB", -- 0x1978
		x"F1",x"FE",x"1F",x"20",x"02",x"3E",x"FF",x"3C", -- 0x1980
		x"E6",x"1C",x"0F",x"4F",x"3A",x"03",x"E1",x"E6", -- 0x1988
		x"03",x"FE",x"03",x"20",x"11",x"21",x"DC",x"98", -- 0x1990
		x"22",x"CE",x"EB",x"21",x"DC",x"98",x"22",x"CA", -- 0x1998
		x"EB",x"21",x"5C",x"97",x"18",x"23",x"21",x"10", -- 0x19A0
		x"80",x"3E",x"02",x"F3",x"32",x"06",x"C8",x"CD", -- 0x19A8
		x"38",x"19",x"22",x"CE",x"EB",x"21",x"00",x"80", -- 0x19B0
		x"CD",x"38",x"19",x"22",x"CA",x"EB",x"21",x"20", -- 0x19B8
		x"80",x"CD",x"38",x"19",x"AF",x"32",x"06",x"C8", -- 0x19C0
		x"FB",x"22",x"C8",x"EB",x"3A",x"03",x"E1",x"4F", -- 0x19C8
		x"2F",x"E6",x"03",x"28",x"0D",x"79",x"E6",x"1C", -- 0x19D0
		x"0F",x"0F",x"4F",x"06",x"00",x"21",x"E0",x"1A", -- 0x19D8
		x"09",x"7E",x"32",x"AF",x"E0",x"3E",x"02",x"32", -- 0x19E0
		x"D5",x"E0",x"3A",x"02",x"E1",x"FE",x"04",x"38", -- 0x19E8
		x"29",x"D6",x"04",x"E6",x"03",x"F5",x"1E",x"00", -- 0x19F0
		x"CB",x"3F",x"30",x"02",x"1E",x"80",x"57",x"3A", -- 0x19F8
		x"AF",x"E0",x"32",x"D5",x"E0",x"2A",x"C8",x"EB", -- 0x1A00
		x"19",x"EB",x"F1",x"FE",x"03",x"20",x"05",x"2A", -- 0x1A08
		x"C8",x"EB",x"18",x"04",x"21",x"80",x"00",x"19", -- 0x1A10
		x"18",x"23",x"11",x"30",x"80",x"21",x"B2",x"80", -- 0x1A18
		x"B7",x"28",x"1A",x"EB",x"21",x"DC",x"98",x"3D", -- 0x1A20
		x"28",x"13",x"08",x"3A",x"AF",x"E0",x"32",x"D5", -- 0x1A28
		x"E0",x"08",x"EB",x"2A",x"CE",x"EB",x"3D",x"28", -- 0x1A30
		x"04",x"EB",x"2A",x"C8",x"EB",x"3E",x"02",x"32", -- 0x1A38
		x"0A",x"E1",x"22",x"D8",x"EB",x"EB",x"22",x"D6", -- 0x1A40
		x"EB",x"3A",x"D5",x"E0",x"32",x"05",x"C8",x"21", -- 0x1A48
		x"48",x"00",x"19",x"22",x"DA",x"EB",x"11",x"00", -- 0x1A50
		x"EA",x"3A",x"D3",x"E0",x"0F",x"30",x"02",x"1E", -- 0x1A58
		x"80",x"2A",x"D6",x"EB",x"01",x"80",x"00",x"3E", -- 0x1A60
		x"02",x"F3",x"32",x"06",x"C8",x"ED",x"B0",x"16", -- 0x1A68
		x"EA",x"2A",x"D8",x"EB",x"01",x"80",x"00",x"3A", -- 0x1A70
		x"0A",x"E1",x"32",x"06",x"C8",x"ED",x"B0",x"AF", -- 0x1A78
		x"32",x"06",x"C8",x"FB",x"21",x"00",x"EA",x"11", -- 0x1A80
		x"00",x"D8",x"3A",x"D3",x"E0",x"0F",x"30",x"06", -- 0x1A88
		x"21",x"80",x"EA",x"11",x"00",x"DA",x"E5",x"D5", -- 0x1A90
		x"CD",x"93",x"0E",x"E1",x"11",x"20",x"00",x"19", -- 0x1A98
		x"EB",x"E1",x"7D",x"C6",x"08",x"E6",x"F8",x"6F", -- 0x1AA0
		x"20",x"EC",x"21",x"C0",x"EA",x"3A",x"D3",x"E0", -- 0x1AA8
		x"0F",x"30",x"03",x"21",x"40",x"EA",x"22",x"C4", -- 0x1AB0
		x"EB",x"2A",x"DA",x"EB",x"22",x"C0",x"EB",x"21", -- 0x1AB8
		x"E1",x"DA",x"3A",x"D3",x"E0",x"0F",x"30",x"03", -- 0x1AC0
		x"21",x"E1",x"D8",x"22",x"C2",x"EB",x"11",x"E0", -- 0x1AC8
		x"EB",x"3A",x"D3",x"E0",x"0F",x"21",x"B8",x"EA", -- 0x1AD0
		x"30",x"03",x"21",x"38",x"EA",x"C3",x"93",x"0E", -- 0x1AD8
		x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"01", -- 0x1AE0
		x"04",x"07",x"2B",x"09",x"34",x"04",x"03",x"B1", -- 0x1AE8
		x"0C",x"04",x"F5",x"2D",x"01",x"AF",x"32",x"99", -- 0x1AF0
		x"E0",x"32",x"98",x"E0",x"32",x"97",x"E0",x"32", -- 0x1AF8
		x"A0",x"E0",x"32",x"A7",x"E0",x"3A",x"02",x"E1", -- 0x1B00
		x"B7",x"28",x"15",x"21",x"80",x"4E",x"22",x"0C", -- 0x1B08
		x"E1",x"3E",x"70",x"32",x"0E",x"E1",x"3E",x"28", -- 0x1B10
		x"32",x"0F",x"E1",x"32",x"FD",x"E0",x"18",x"06", -- 0x1B18
		x"21",x"B7",x"0E",x"22",x"0C",x"E1",x"DD",x"21", -- 0x1B20
		x"20",x"E1",x"DD",x"CB",x"00",x"EE",x"AF",x"DD", -- 0x1B28
		x"77",x"06",x"DD",x"21",x"30",x"E1",x"DD",x"CB", -- 0x1B30
		x"00",x"EE",x"DD",x"77",x"06",x"3A",x"02",x"E1", -- 0x1B38
		x"B7",x"20",x"7E",x"3E",x"01",x"32",x"98",x"E0", -- 0x1B40
		x"32",x"93",x"E0",x"3A",x"00",x"E1",x"CB",x"6F", -- 0x1B48
		x"28",x"08",x"06",x"02",x"DF",x"CD",x"AE",x"20", -- 0x1B50
		x"30",x"F8",x"3A",x"00",x"E1",x"CB",x"6F",x"20", -- 0x1B58
		x"0A",x"3E",x"78",x"32",x"0E",x"E1",x"3E",x"28", -- 0x1B60
		x"32",x"0F",x"E1",x"3E",x"31",x"32",x"FD",x"E0", -- 0x1B68
		x"3E",x"02",x"01",x"BB",x"20",x"FF",x"3E",x"0E", -- 0x1B70
		x"01",x"82",x"17",x"FF",x"0E",x"0D",x"CD",x"78", -- 0x1B78
		x"11",x"21",x"75",x"1E",x"CD",x"DF",x"1C",x"CD", -- 0x1B80
		x"3A",x"29",x"06",x"01",x"DF",x"CD",x"4A",x"1D", -- 0x1B88
		x"CD",x"3A",x"29",x"06",x"01",x"DF",x"3A",x"93", -- 0x1B90
		x"E0",x"B7",x"20",x"F1",x"32",x"98",x"E0",x"0E", -- 0x1B98
		x"06",x"CD",x"78",x"11",x"CD",x"02",x"1D",x"21", -- 0x1BA0
		x"B5",x"1E",x"CD",x"DF",x"1C",x"CD",x"4A",x"1D", -- 0x1BA8
		x"CD",x"BA",x"1C",x"CD",x"3A",x"29",x"06",x"01", -- 0x1BB0
		x"DF",x"3A",x"93",x"E0",x"B7",x"20",x"EE",x"18", -- 0x1BB8
		x"1B",x"3E",x"02",x"01",x"BB",x"20",x"FF",x"3E", -- 0x1BC0
		x"0E",x"01",x"82",x"17",x"FF",x"3A",x"03",x"E1", -- 0x1BC8
		x"2F",x"E6",x"03",x"0E",x"12",x"20",x"02",x"0E", -- 0x1BD0
		x"13",x"CD",x"78",x"11",x"AF",x"32",x"C5",x"E0", -- 0x1BD8
		x"0E",x"0C",x"CD",x"78",x"11",x"06",x"01",x"DF", -- 0x1BE0
		x"CD",x"BA",x"1C",x"3A",x"26",x"E1",x"B7",x"28", -- 0x1BE8
		x"F4",x"3A",x"36",x"E1",x"B7",x"28",x"EE",x"AF", -- 0x1BF0
		x"32",x"A7",x"E0",x"CD",x"35",x"2D",x"32",x"A0", -- 0x1BF8
		x"E0",x"4F",x"3A",x"F0",x"E0",x"81",x"32",x"F0", -- 0x1C00
		x"E0",x"3A",x"93",x"E0",x"0F",x"DA",x"3C",x"1D", -- 0x1C08
		x"3A",x"99",x"E0",x"B7",x"C2",x"7F",x"1F",x"3A", -- 0x1C10
		x"A0",x"E0",x"E6",x"20",x"28",x"0E",x"21",x"9B", -- 0x1C18
		x"E0",x"7E",x"B7",x"28",x"07",x"35",x"CD",x"67", -- 0x1C20
		x"18",x"C3",x"CA",x"1C",x"CD",x"96",x"25",x"3A", -- 0x1C28
		x"A9",x"E0",x"B7",x"C4",x"BE",x"1F",x"CD",x"17", -- 0x1C30
		x"27",x"3A",x"18",x"E1",x"E6",x"03",x"C4",x"E8", -- 0x1C38
		x"28",x"CD",x"BA",x"1C",x"3A",x"99",x"E0",x"FE", -- 0x1C40
		x"03",x"D2",x"9D",x"1C",x"3A",x"93",x"E0",x"B7", -- 0x1C48
		x"28",x"08",x"3A",x"97",x"E0",x"FE",x"0F",x"DA", -- 0x1C50
		x"9D",x"1C",x"3A",x"A1",x"E0",x"FE",x"03",x"D2", -- 0x1C58
		x"9D",x"1C",x"3A",x"A0",x"E0",x"E6",x"10",x"20", -- 0x1C60
		x"06",x"32",x"A2",x"E0",x"C3",x"9D",x"1C",x"21", -- 0x1C68
		x"F0",x"E0",x"34",x"21",x"A3",x"E0",x"3A",x"A2", -- 0x1C70
		x"E0",x"E6",x"01",x"28",x"17",x"34",x"7E",x"3D", -- 0x1C78
		x"28",x"08",x"FE",x"41",x"30",x"15",x"FE",x"20", -- 0x1C80
		x"20",x"13",x"CD",x"46",x"29",x"0E",x"05",x"CD", -- 0x1C88
		x"78",x"11",x"18",x"09",x"77",x"3C",x"32",x"A2", -- 0x1C90
		x"E0",x"18",x"02",x"36",x"1F",x"DD",x"21",x"60", -- 0x1C98
		x"E2",x"06",x"03",x"C5",x"DD",x"7E",x"00",x"CB", -- 0x1CA0
		x"47",x"C2",x"1C",x"2A",x"01",x"10",x"00",x"DD", -- 0x1CA8
		x"09",x"C1",x"10",x"EF",x"06",x"01",x"DF",x"C3", -- 0x1CB0
		x"F7",x"1B",x"21",x"AD",x"E0",x"35",x"C0",x"36", -- 0x1CB8
		x"02",x"3A",x"0D",x"E1",x"EE",x"01",x"32",x"0D", -- 0x1CC0
		x"E1",x"C9",x"AF",x"32",x"A1",x"E0",x"0E",x"06", -- 0x1CC8
		x"CD",x"78",x"11",x"CD",x"D9",x"1C",x"C3",x"2F", -- 0x1CD0
		x"1C",x"CD",x"02",x"1D",x"21",x"1E",x"1F",x"AF", -- 0x1CD8
		x"32",x"97",x"E0",x"CD",x"8A",x"1D",x"21",x"A5", -- 0x1CE0
		x"E0",x"CB",x"CE",x"3A",x"98",x"E0",x"B7",x"C0", -- 0x1CE8
		x"3A",x"99",x"E0",x"B7",x"CA",x"C1",x"25",x"3A", -- 0x1CF0
		x"A7",x"E0",x"E6",x"0C",x"32",x"A7",x"E0",x"C3", -- 0x1CF8
		x"C1",x"25",x"AF",x"32",x"60",x"E2",x"32",x"70", -- 0x1D00
		x"E2",x"32",x"80",x"E2",x"67",x"6F",x"22",x"05", -- 0x1D08
		x"EB",x"22",x"09",x"EB",x"22",x"0D",x"EB",x"21", -- 0x1D10
		x"93",x"E0",x"CB",x"C6",x"3A",x"B4",x"E7",x"B7", -- 0x1D18
		x"C0",x"21",x"48",x"EB",x"11",x"49",x"EB",x"36", -- 0x1D20
		x"00",x"01",x"18",x"00",x"ED",x"B0",x"21",x"68", -- 0x1D28
		x"EB",x"11",x"69",x"EB",x"36",x"00",x"01",x"18", -- 0x1D30
		x"00",x"ED",x"B0",x"C9",x"3A",x"99",x"E0",x"FE", -- 0x1D38
		x"01",x"CC",x"94",x"1F",x"CD",x"4A",x"1D",x"C3", -- 0x1D40
		x"2F",x"1C",x"2A",x"94",x"E0",x"ED",x"4B",x"7C", -- 0x1D48
		x"E1",x"09",x"5C",x"26",x"00",x"22",x"7C",x"E1", -- 0x1D50
		x"3A",x"96",x"E0",x"B7",x"3A",x"0F",x"E1",x"C2", -- 0x1D58
		x"66",x"1D",x"83",x"C3",x"67",x"1D",x"93",x"32", -- 0x1D60
		x"0F",x"E1",x"21",x"92",x"E0",x"35",x"20",x"17", -- 0x1D68
		x"2A",x"90",x"E0",x"CD",x"8A",x"1D",x"30",x"0F", -- 0x1D70
		x"21",x"93",x"E0",x"CB",x"86",x"21",x"99",x"E0", -- 0x1D78
		x"7E",x"FE",x"04",x"C2",x"87",x"1D",x"34",x"C3", -- 0x1D80
		x"EB",x"1C",x"7E",x"B7",x"CA",x"2C",x"1E",x"FE", -- 0x1D88
		x"FF",x"CA",x"33",x"1E",x"5F",x"E6",x"3F",x"32", -- 0x1D90
		x"92",x"E0",x"CB",x"7B",x"CA",x"09",x"1E",x"23", -- 0x1D98
		x"7E",x"32",x"0C",x"E1",x"47",x"23",x"7E",x"32", -- 0x1DA0
		x"0D",x"E1",x"4F",x"23",x"3A",x"97",x"E0",x"3C", -- 0x1DA8
		x"32",x"97",x"E0",x"CB",x"5E",x"28",x"0F",x"CB", -- 0x1DB0
		x"56",x"16",x"08",x"28",x"02",x"16",x"F8",x"3A", -- 0x1DB8
		x"0E",x"E1",x"82",x"32",x"0E",x"E1",x"CB",x"4E", -- 0x1DC0
		x"28",x"0F",x"CB",x"46",x"16",x"08",x"28",x"02", -- 0x1DC8
		x"16",x"F8",x"3A",x"0F",x"E1",x"82",x"32",x"0F", -- 0x1DD0
		x"E1",x"3A",x"99",x"E0",x"FE",x"03",x"30",x"29", -- 0x1DD8
		x"B7",x"20",x"06",x"3A",x"98",x"E0",x"B7",x"20", -- 0x1DE0
		x"20",x"3A",x"97",x"E0",x"FE",x"06",x"38",x"19", -- 0x1DE8
		x"FE",x"0B",x"20",x"09",x"AF",x"32",x"05",x"EB", -- 0x1DF0
		x"32",x"06",x"EB",x"18",x"0C",x"30",x"0A",x"78", -- 0x1DF8
		x"D6",x"08",x"32",x"04",x"EB",x"79",x"32",x"05", -- 0x1E00
		x"EB",x"23",x"4E",x"23",x"46",x"23",x"22",x"90", -- 0x1E08
		x"E0",x"ED",x"43",x"94",x"E0",x"3A",x"96",x"E0", -- 0x1E10
		x"57",x"7B",x"E6",x"40",x"BA",x"CA",x"2A",x"1E", -- 0x1E18
		x"32",x"96",x"E0",x"AF",x"32",x"7C",x"E1",x"32", -- 0x1E20
		x"7D",x"E1",x"B7",x"C9",x"21",x"A5",x"E0",x"CB", -- 0x1E28
		x"8E",x"37",x"C9",x"23",x"3A",x"0F",x"E1",x"BE", -- 0x1E30
		x"23",x"DA",x"8A",x"1D",x"3E",x"01",x"32",x"92", -- 0x1E38
		x"E0",x"C3",x"2A",x"1E",x"8A",x"A6",x"4E",x"00", -- 0x1E40
		x"00",x"00",x"8A",x"AE",x"4E",x"00",x"00",x"00", -- 0x1E48
		x"8C",x"F8",x"4E",x"00",x"00",x"00",x"8E",x"B6", -- 0x1E50
		x"0E",x"08",x"00",x"00",x"01",x"00",x"00",x"01", -- 0x1E58
		x"00",x"00",x"90",x"B7",x"0E",x"00",x"00",x"00", -- 0x1E60
		x"1E",x"80",x"00",x"1E",x"40",x"00",x"1E",x"20", -- 0x1E68
		x"00",x"02",x"00",x"00",x"00",x"90",x"B7",x"0E", -- 0x1E70
		x"00",x"40",x"00",x"90",x"B7",x"0E",x"00",x"40", -- 0x1E78
		x"00",x"0A",x"40",x"00",x"0A",x"80",x"00",x"10", -- 0x1E80
		x"C0",x"00",x"8E",x"B7",x"0E",x"00",x"C0",x"00", -- 0x1E88
		x"84",x"B6",x"0E",x"00",x"C0",x"00",x"84",x"F8", -- 0x1E90
		x"4E",x"0C",x"00",x"01",x"84",x"AE",x"4E",x"00", -- 0x1E98
		x"00",x"01",x"84",x"A6",x"4E",x"00",x"40",x"01", -- 0x1EA0
		x"84",x"80",x"4E",x"00",x"80",x"01",x"84",x"80", -- 0x1EA8
		x"4E",x"00",x"80",x"01",x"00",x"88",x"90",x"4E", -- 0x1EB0
		x"00",x"C0",x"00",x"88",x"98",x"4E",x"00",x"80", -- 0x1EB8
		x"00",x"C8",x"92",x"4E",x"00",x"50",x"00",x"C8", -- 0x1EC0
		x"9A",x"4E",x"00",x"00",x"00",x"C7",x"94",x"4E", -- 0x1EC8
		x"00",x"50",x"00",x"C7",x"AA",x"4E",x"03",x"80", -- 0x1ED0
		x"00",x"C7",x"AC",x"4E",x"00",x"C0",x"00",x"C8", -- 0x1ED8
		x"C8",x"4E",x"00",x"00",x"01",x"48",x"80",x"01", -- 0x1EE0
		x"FF",x"28",x"48",x"00",x"01",x"C8",x"CA",x"4E", -- 0x1EE8
		x"00",x"C0",x"00",x"C8",x"CC",x"4E",x"00",x"80", -- 0x1EF0
		x"00",x"C8",x"9C",x"4E",x"02",x"50",x"00",x"C8", -- 0x1EF8
		x"96",x"4E",x"00",x"00",x"00",x"88",x"9E",x"4E", -- 0x1F00
		x"00",x"50",x"00",x"88",x"A0",x"4E",x"00",x"80", -- 0x1F08
		x"00",x"8A",x"A8",x"4E",x"00",x"C0",x"00",x"88", -- 0x1F10
		x"80",x"4E",x"00",x"00",x"01",x"00",x"88",x"90", -- 0x1F18
		x"4E",x"00",x"C0",x"00",x"88",x"98",x"4E",x"00", -- 0x1F20
		x"80",x"00",x"C8",x"92",x"4E",x"00",x"50",x"00", -- 0x1F28
		x"C8",x"9A",x"4E",x"00",x"00",x"00",x"C7",x"94", -- 0x1F30
		x"4E",x"00",x"50",x"00",x"C7",x"AA",x"4E",x"03", -- 0x1F38
		x"80",x"00",x"C7",x"AC",x"4E",x"00",x"C0",x"00", -- 0x1F40
		x"C8",x"C8",x"4E",x"00",x"00",x"01",x"C7",x"CA", -- 0x1F48
		x"4E",x"00",x"C0",x"00",x"C7",x"CC",x"4E",x"00", -- 0x1F50
		x"80",x"00",x"C8",x"9C",x"4E",x"02",x"50",x"00", -- 0x1F58
		x"C8",x"96",x"4E",x"00",x"00",x"00",x"88",x"9E", -- 0x1F60
		x"4E",x"00",x"50",x"00",x"88",x"A0",x"4E",x"00", -- 0x1F68
		x"80",x"00",x"8A",x"A8",x"4E",x"00",x"C0",x"00", -- 0x1F70
		x"88",x"80",x"4E",x"00",x"00",x"01",x"00",x"3D", -- 0x1F78
		x"E6",x"07",x"CD",x"F7",x"66",x"8F",x"1F",x"E7", -- 0x1F80
		x"1F",x"22",x"20",x"58",x"20",x"61",x"20",x"CD", -- 0x1F88
		x"94",x"1F",x"18",x"53",x"3E",x"01",x"32",x"A5", -- 0x1F90
		x"E0",x"0E",x"10",x"CD",x"78",x"11",x"DD",x"21", -- 0x1F98
		x"58",x"A2",x"CD",x"CC",x"2C",x"21",x"41",x"D0", -- 0x1FA0
		x"01",x"1D",x"1C",x"16",x"30",x"CD",x"53",x"02", -- 0x1FA8
		x"CD",x"C6",x"1F",x"3E",x"05",x"01",x"5C",x"22", -- 0x1FB0
		x"FF",x"21",x"99",x"E0",x"34",x"C9",x"CB",x"7F", -- 0x1FB8
		x"C0",x"CB",x"FF",x"32",x"A9",x"E0",x"AF",x"32", -- 0x1FC0
		x"A6",x"E9",x"DD",x"21",x"20",x"E1",x"DD",x"77", -- 0x1FC8
		x"06",x"DD",x"CB",x"00",x"E6",x"DD",x"21",x"30", -- 0x1FD0
		x"E1",x"DD",x"77",x"06",x"DD",x"CB",x"00",x"E6", -- 0x1FD8
		x"3E",x"02",x"01",x"9B",x"21",x"FF",x"C9",x"0E", -- 0x1FE0
		x"00",x"2A",x"0E",x"E1",x"7D",x"E6",x"FE",x"FE", -- 0x1FE8
		x"70",x"28",x"06",x"0E",x"02",x"30",x"02",x"0E", -- 0x1FF0
		x"01",x"7C",x"FE",x"60",x"30",x"0B",x"E6",x"FE", -- 0x1FF8
		x"FE",x"5E",x"CA",x"09",x"20",x"3E",x"08",x"B1", -- 0x2000
		x"4F",x"21",x"9A",x"E0",x"7E",x"B7",x"28",x"04", -- 0x2008
		x"35",x"AF",x"18",x"08",x"79",x"B7",x"20",x"04", -- 0x2010
		x"21",x"99",x"E0",x"34",x"32",x"A0",x"E0",x"C3", -- 0x2018
		x"2C",x"1C",x"3A",x"02",x"E1",x"B7",x"28",x"0F", -- 0x2020
		x"FE",x"44",x"30",x"0B",x"FE",x"43",x"38",x"22", -- 0x2028
		x"3A",x"D2",x"E0",x"FE",x"40",x"38",x"1B",x"21", -- 0x2030
		x"99",x"E0",x"34",x"AF",x"32",x"97",x"E0",x"32", -- 0x2038
		x"A0",x"E0",x"21",x"93",x"E0",x"CB",x"CE",x"0E", -- 0x2040
		x"0F",x"CD",x"78",x"11",x"21",x"44",x"1E",x"CD", -- 0x2048
		x"DF",x"1C",x"CD",x"3A",x"29",x"C3",x"41",x"1C", -- 0x2050
		x"AF",x"32",x"A0",x"E0",x"CD",x"4A",x"1D",x"18", -- 0x2058
		x"F1",x"06",x"01",x"DF",x"3A",x"A6",x"E9",x"E6", -- 0x2060
		x"03",x"FE",x"03",x"20",x"F4",x"0E",x"10",x"CD", -- 0x2068
		x"78",x"11",x"0E",x"00",x"CD",x"78",x"11",x"06", -- 0x2070
		x"02",x"DF",x"CD",x"AE",x"20",x"3A",x"A6",x"E9", -- 0x2078
		x"07",x"30",x"F4",x"21",x"41",x"D0",x"01",x"1D", -- 0x2080
		x"1C",x"16",x"30",x"CD",x"53",x"02",x"AF",x"32", -- 0x2088
		x"13",x"E1",x"21",x"10",x"EB",x"11",x"11",x"EB", -- 0x2090
		x"01",x"6F",x"00",x"77",x"ED",x"B0",x"21",x"00", -- 0x2098
		x"E1",x"CB",x"EE",x"3A",x"03",x"E1",x"FE",x"20", -- 0x20A0
		x"DA",x"FE",x"14",x"C3",x"F7",x"6F",x"21",x"0F", -- 0x20A8
		x"E1",x"7E",x"FE",x"81",x"D8",x"35",x"CD",x"3A", -- 0x20B0
		x"29",x"B7",x"C9",x"CD",x"32",x"22",x"DA",x"EE", -- 0x20B8
		x"20",x"DD",x"21",x"20",x"E1",x"CD",x"1A",x"21", -- 0x20C0
		x"DD",x"21",x"30",x"E1",x"CD",x"1A",x"21",x"06", -- 0x20C8
		x"01",x"DF",x"DD",x"21",x"20",x"E1",x"CD",x"3D", -- 0x20D0
		x"21",x"DD",x"21",x"30",x"E1",x"CD",x"3D",x"21", -- 0x20D8
		x"DD",x"7E",x"06",x"E6",x"01",x"28",x"E8",x"3A", -- 0x20E0
		x"26",x"E1",x"E6",x"01",x"28",x"E1",x"3A",x"C5", -- 0x20E8
		x"E0",x"B7",x"28",x"1B",x"DD",x"21",x"20",x"E1", -- 0x20F0
		x"DD",x"CB",x"00",x"7E",x"C4",x"55",x"27",x"DD", -- 0x20F8
		x"21",x"30",x"E1",x"DD",x"CB",x"00",x"7E",x"C4", -- 0x2100
		x"55",x"27",x"06",x"01",x"DF",x"18",x"DF",x"21", -- 0x2108
		x"20",x"E1",x"CB",x"AE",x"21",x"30",x"E1",x"CB", -- 0x2110
		x"AE",x"F7",x"DD",x"CB",x"00",x"7E",x"C8",x"DD", -- 0x2118
		x"36",x"0C",x"00",x"DD",x"36",x"0D",x"12",x"DD", -- 0x2120
		x"36",x"0F",x"F1",x"DD",x"CB",x"00",x"76",x"3E", -- 0x2128
		x"63",x"28",x"02",x"3E",x"8D",x"DD",x"77",x"0E", -- 0x2130
		x"DD",x"36",x"05",x"02",x"C9",x"DD",x"CB",x"00", -- 0x2138
		x"7E",x"C8",x"3A",x"FD",x"E0",x"57",x"3A",x"02", -- 0x2140
		x"E1",x"B7",x"28",x"04",x"3A",x"0F",x"E1",x"57", -- 0x2148
		x"DD",x"CB",x"0D",x"66",x"20",x"1E",x"DD",x"7E", -- 0x2150
		x"0F",x"BA",x"30",x"35",x"01",x"C0",x"00",x"C6", -- 0x2158
		x"08",x"BA",x"30",x"13",x"C6",x"08",x"01",x"00", -- 0x2160
		x"01",x"BA",x"30",x"0B",x"C6",x"08",x"01",x"80", -- 0x2168
		x"01",x"BA",x"30",x"03",x"01",x"00",x"02",x"3A", -- 0x2170
		x"FC",x"E0",x"6F",x"26",x"00",x"09",x"7D",x"32", -- 0x2178
		x"FC",x"E0",x"DD",x"7E",x"0F",x"84",x"DD",x"77", -- 0x2180
		x"0F",x"30",x"0D",x"DD",x"CB",x"0D",x"A6",x"18", -- 0x2188
		x"07",x"DD",x"72",x"0F",x"DD",x"CB",x"06",x"C6", -- 0x2190
		x"C3",x"55",x"27",x"CD",x"32",x"22",x"DA",x"D3", -- 0x2198
		x"21",x"21",x"66",x"87",x"CD",x"24",x"22",x"06", -- 0x21A0
		x"01",x"DF",x"DD",x"21",x"20",x"E1",x"CD",x"D9", -- 0x21A8
		x"21",x"DD",x"21",x"30",x"E1",x"CD",x"D9",x"21", -- 0x21B0
		x"21",x"FB",x"E0",x"35",x"20",x"07",x"2A",x"F8", -- 0x21B8
		x"E0",x"23",x"CD",x"24",x"22",x"DD",x"7E",x"06", -- 0x21C0
		x"E6",x"01",x"28",x"DB",x"3A",x"26",x"E1",x"E6", -- 0x21C8
		x"01",x"28",x"D4",x"21",x"A6",x"E9",x"CB",x"CE", -- 0x21D0
		x"F7",x"DD",x"CB",x"06",x"46",x"C0",x"2A",x"F8", -- 0x21D8
		x"E0",x"5E",x"16",x"00",x"42",x"EB",x"29",x"29", -- 0x21E0
		x"3A",x"FC",x"E0",x"4F",x"09",x"EB",x"7B",x"32", -- 0x21E8
		x"FC",x"E0",x"DD",x"7E",x"0F",x"CB",x"46",x"20", -- 0x21F0
		x"03",x"82",x"18",x"01",x"92",x"DD",x"77",x"0F", -- 0x21F8
		x"30",x"04",x"DD",x"CB",x"0D",x"E6",x"DD",x"CB", -- 0x2200
		x"0D",x"66",x"28",x"0F",x"FE",x"F1",x"30",x"0B", -- 0x2208
		x"DD",x"CB",x"06",x"C6",x"AF",x"DD",x"77",x"0E", -- 0x2210
		x"DD",x"77",x"0E",x"3A",x"FA",x"E0",x"DD",x"77", -- 0x2218
		x"0C",x"C3",x"55",x"27",x"7E",x"32",x"FB",x"E0", -- 0x2220
		x"23",x"7E",x"32",x"FA",x"E0",x"23",x"22",x"F8", -- 0x2228
		x"E0",x"C9",x"16",x"00",x"DD",x"21",x"20",x"E1", -- 0x2230
		x"DD",x"7E",x"00",x"E6",x"8E",x"FE",x"82",x"28", -- 0x2238
		x"05",x"DD",x"CB",x"06",x"C6",x"14",x"DD",x"21", -- 0x2240
		x"30",x"E1",x"DD",x"7E",x"00",x"E6",x"8E",x"FE", -- 0x2248
		x"82",x"28",x"07",x"DD",x"CB",x"06",x"C6",x"7A", -- 0x2250
		x"0F",x"C9",x"B7",x"C9",x"3A",x"03",x"E1",x"2F", -- 0x2258
		x"E6",x"03",x"0E",x"15",x"CC",x"78",x"11",x"CD", -- 0x2260
		x"88",x"25",x"CD",x"64",x"24",x"21",x"65",x"E1", -- 0x2268
		x"11",x"6C",x"E7",x"01",x"03",x"00",x"ED",x"B0", -- 0x2270
		x"CD",x"C1",x"24",x"3A",x"74",x"E7",x"32",x"7F", -- 0x2278
		x"E7",x"21",x"78",x"E7",x"CD",x"BE",x"23",x"CD", -- 0x2280
		x"F2",x"23",x"21",x"D1",x"A5",x"CD",x"70",x"23", -- 0x2288
		x"21",x"B4",x"D2",x"11",x"78",x"E7",x"06",x"03", -- 0x2290
		x"CD",x"96",x"23",x"06",x"01",x"3E",x"29",x"CD", -- 0x2298
		x"B1",x"23",x"06",x"0A",x"DF",x"0E",x"1B",x"CD", -- 0x22A0
		x"78",x"11",x"21",x"68",x"E7",x"01",x"08",x"00", -- 0x22A8
		x"50",x"CD",x"E2",x"01",x"21",x"02",x"A6",x"3A", -- 0x22B0
		x"7F",x"E7",x"FE",x"32",x"38",x"65",x"21",x"0E", -- 0x22B8
		x"A6",x"FE",x"64",x"30",x"4B",x"D6",x"32",x"0E", -- 0x22C0
		x"00",x"FE",x"05",x"38",x"05",x"D6",x"05",x"0C", -- 0x22C8
		x"18",x"F7",x"CB",x"01",x"06",x"00",x"21",x"5C", -- 0x22D0
		x"23",x"09",x"11",x"6B",x"E7",x"DD",x"21",x"8C", -- 0x22D8
		x"D1",x"06",x"02",x"7E",x"DD",x"77",x"00",x"FE", -- 0x22E0
		x"30",x"20",x"01",x"AF",x"12",x"13",x"23",x"C5", -- 0x22E8
		x"01",x"20",x"00",x"DD",x"09",x"C1",x"10",x"EB", -- 0x22F0
		x"21",x"CE",x"D1",x"11",x"1A",x"A6",x"06",x"05", -- 0x22F8
		x"CD",x"EE",x"01",x"21",x"CC",x"D1",x"11",x"24", -- 0x2300
		x"A6",x"06",x"07",x"CD",x"EE",x"01",x"18",x"08", -- 0x2308
		x"CD",x"22",x"02",x"3E",x"05",x"32",x"6B",x"E7", -- 0x2310
		x"21",x"6F",x"E7",x"CD",x"D1",x"12",x"CD",x"55", -- 0x2318
		x"2D",x"18",x"03",x"CD",x"22",x"02",x"3A",x"9B", -- 0x2320
		x"E0",x"B7",x"28",x"27",x"32",x"6C",x"E7",x"AF", -- 0x2328
		x"32",x"6B",x"E7",x"21",x"66",x"A6",x"CD",x"22", -- 0x2330
		x"02",x"3A",x"6C",x"E7",x"32",x"09",x"D2",x"21", -- 0x2338
		x"29",x"D2",x"11",x"24",x"A6",x"06",x"07",x"CD", -- 0x2340
		x"EE",x"01",x"21",x"6F",x"E7",x"CD",x"D1",x"12", -- 0x2348
		x"CD",x"55",x"2D",x"06",x"3C",x"DF",x"21",x"A6", -- 0x2350
		x"E9",x"CB",x"C6",x"F7",x"30",x"01",x"30",x"01", -- 0x2358
		x"30",x"02",x"30",x"02",x"30",x"03",x"30",x"03", -- 0x2360
		x"30",x"04",x"30",x"05",x"01",x"00",x"02",x"00", -- 0x2368
		x"46",x"23",x"4E",x"AF",x"B9",x"C8",x"23",x"5E", -- 0x2370
		x"23",x"56",x"23",x"EB",x"C5",x"DF",x"1A",x"FE", -- 0x2378
		x"30",x"F5",x"06",x"01",x"CD",x"EE",x"01",x"F1", -- 0x2380
		x"0E",x"09",x"E5",x"C4",x"78",x"11",x"E1",x"C1", -- 0x2388
		x"0D",x"20",x"E9",x"EB",x"18",x"DC",x"C5",x"1A", -- 0x2390
		x"FE",x"30",x"F5",x"28",x"03",x"06",x"0A",x"DF", -- 0x2398
		x"06",x"01",x"CD",x"EE",x"01",x"F1",x"0E",x"09", -- 0x23A0
		x"E5",x"C4",x"78",x"11",x"E1",x"C1",x"10",x"E6", -- 0x23A8
		x"C9",x"F5",x"06",x"0A",x"DF",x"F1",x"CD",x"EA", -- 0x23B0
		x"01",x"0E",x"09",x"C3",x"78",x"11",x"01",x"00", -- 0x23B8
		x"01",x"51",x"FE",x"64",x"30",x"0B",x"05",x"FE", -- 0x23C0
		x"0A",x"38",x"05",x"D6",x"0A",x"0C",x"18",x"F7", -- 0x23C8
		x"57",x"1E",x"00",x"78",x"CD",x"DD",x"23",x"79", -- 0x23D0
		x"CD",x"DD",x"23",x"72",x"C9",x"B7",x"20",x"09", -- 0x23D8
		x"CB",x"43",x"20",x"02",x"3E",x"30",x"77",x"23", -- 0x23E0
		x"C9",x"CB",x"C3",x"18",x"F9",x"21",x"4D",x"E1", -- 0x23E8
		x"18",x"03",x"21",x"55",x"E1",x"11",x"68",x"E7", -- 0x23F0
		x"01",x"03",x"00",x"ED",x"B0",x"21",x"60",x"E7", -- 0x23F8
		x"11",x"61",x"E7",x"01",x"07",x"00",x"36",x"00", -- 0x2400
		x"ED",x"B0",x"FD",x"21",x"4F",x"24",x"06",x"07", -- 0x2408
		x"11",x"60",x"E7",x"C5",x"2A",x"68",x"E7",x"3A", -- 0x2410
		x"6A",x"E7",x"FD",x"4E",x"00",x"FD",x"46",x"01", -- 0x2418
		x"B7",x"ED",x"42",x"FD",x"9E",x"02",x"38",x"0B", -- 0x2420
		x"22",x"68",x"E7",x"32",x"6A",x"E7",x"EB",x"34", -- 0x2428
		x"EB",x"18",x"ED",x"FD",x"23",x"FD",x"23",x"FD", -- 0x2430
		x"23",x"13",x"C1",x"10",x"D6",x"3A",x"68",x"E7", -- 0x2438
		x"12",x"21",x"60",x"E7",x"1E",x"00",x"06",x"07", -- 0x2440
		x"7E",x"CD",x"DD",x"23",x"10",x"FA",x"C9",x"80", -- 0x2448
		x"96",x"98",x"40",x"42",x"0F",x"A0",x"86",x"01", -- 0x2450
		x"10",x"27",x"00",x"E8",x"03",x"00",x"64",x"00", -- 0x2458
		x"00",x"0A",x"00",x"00",x"2A",x"55",x"E1",x"3A", -- 0x2460
		x"57",x"E1",x"18",x"06",x"2A",x"4D",x"E1",x"3A", -- 0x2468
		x"4F",x"E1",x"5F",x"AF",x"57",x"06",x"02",x"CD", -- 0x2470
		x"B9",x"24",x"22",x"78",x"E7",x"ED",x"53",x"7A", -- 0x2478
		x"E7",x"06",x"03",x"CD",x"B9",x"24",x"22",x"7C", -- 0x2480
		x"E7",x"ED",x"53",x"7E",x"E7",x"29",x"EB",x"ED", -- 0x2488
		x"6A",x"EB",x"ED",x"4B",x"78",x"E7",x"09",x"22", -- 0x2490
		x"78",x"E7",x"ED",x"4B",x"7A",x"E7",x"EB",x"ED", -- 0x2498
		x"4A",x"22",x"7A",x"E7",x"EB",x"ED",x"4B",x"7C", -- 0x24A0
		x"E7",x"09",x"22",x"64",x"E7",x"ED",x"4B",x"7E", -- 0x24A8
		x"E7",x"EB",x"ED",x"4A",x"22",x"66",x"E7",x"EB", -- 0x24B0
		x"C9",x"29",x"EB",x"ED",x"6A",x"EB",x"10",x"F9", -- 0x24B8
		x"C9",x"CD",x"0B",x"25",x"3E",x"40",x"92",x"47", -- 0x24C0
		x"C5",x"CD",x"E9",x"24",x"38",x"0C",x"C5",x"CD", -- 0x24C8
		x"FA",x"24",x"CD",x"77",x"25",x"C1",x"78",x"B7", -- 0x24D0
		x"28",x"0D",x"CD",x"5F",x"25",x"21",x"6F",x"E7", -- 0x24D8
		x"CD",x"62",x"25",x"C1",x"10",x"E2",x"C9",x"C1", -- 0x24E0
		x"C9",x"06",x"08",x"21",x"6F",x"E7",x"11",x"67", -- 0x24E8
		x"E7",x"1A",x"BE",x"D8",x"C0",x"1B",x"2B",x"10", -- 0x24F0
		x"F8",x"D0",x"06",x"08",x"21",x"68",x"E7",x"11", -- 0x24F8
		x"60",x"E7",x"AF",x"1A",x"9E",x"12",x"13",x"23", -- 0x2500
		x"10",x"F9",x"C9",x"21",x"78",x"E7",x"11",x"79", -- 0x2508
		x"E7",x"36",x"00",x"01",x"07",x"00",x"ED",x"B0", -- 0x2510
		x"3E",x"01",x"32",x"7C",x"E7",x"21",x"67",x"E7", -- 0x2518
		x"CD",x"4E",x"25",x"53",x"21",x"6F",x"E7",x"CD", -- 0x2520
		x"4E",x"25",x"7B",x"BA",x"C8",x"38",x"0F",x"92", -- 0x2528
		x"5F",x"CD",x"6B",x"25",x"21",x"68",x"E7",x"CD", -- 0x2530
		x"6E",x"25",x"1D",x"20",x"F4",x"C9",x"7A",x"93", -- 0x2538
		x"5F",x"CD",x"5F",x"25",x"21",x"6F",x"E7",x"CD", -- 0x2540
		x"62",x"25",x"1D",x"20",x"F4",x"C9",x"0E",x"04", -- 0x2548
		x"1E",x"01",x"06",x"08",x"7E",x"07",x"D8",x"1C", -- 0x2550
		x"10",x"FB",x"2B",x"0D",x"20",x"F4",x"C9",x"21", -- 0x2558
		x"7F",x"E7",x"06",x"08",x"AF",x"CB",x"1E",x"2B", -- 0x2560
		x"10",x"FB",x"C9",x"21",x"78",x"E7",x"06",x"08", -- 0x2568
		x"AF",x"CB",x"16",x"23",x"10",x"FB",x"C9",x"21", -- 0x2570
		x"78",x"E7",x"11",x"70",x"E7",x"06",x"08",x"AF", -- 0x2578
		x"1A",x"8E",x"12",x"23",x"13",x"10",x"F9",x"C9", -- 0x2580
		x"21",x"60",x"E7",x"11",x"61",x"E7",x"01",x"17", -- 0x2588
		x"00",x"36",x"00",x"ED",x"B0",x"C9",x"0E",x"08", -- 0x2590
		x"3A",x"A0",x"E0",x"E6",x"0C",x"28",x"13",x"E6", -- 0x2598
		x"08",x"3A",x"0F",x"E1",x"28",x"08",x"FE",x"A0", -- 0x25A0
		x"30",x"08",x"0E",x"08",x"18",x"0F",x"FE",x"1D", -- 0x25A8
		x"30",x"09",x"AF",x"32",x"7C",x"E1",x"32",x"7D", -- 0x25B0
		x"E1",x"18",x"06",x"0E",x"04",x"79",x"32",x"A7", -- 0x25B8
		x"E0",x"3A",x"A0",x"E0",x"E6",x"03",x"20",x"0A", -- 0x25C0
		x"AF",x"32",x"7E",x"E1",x"32",x"7F",x"E1",x"C3", -- 0x25C8
		x"17",x"26",x"E6",x"02",x"28",x"1E",x"3A",x"20", -- 0x25D0
		x"E1",x"B7",x"06",x"0E",x"28",x"0C",x"CB",x"67", -- 0x25D8
		x"28",x"06",x"3A",x"26",x"E1",x"B7",x"20",x"02", -- 0x25E0
		x"06",x"1E",x"3A",x"0E",x"E1",x"B8",x"38",x"D8", -- 0x25E8
		x"0E",x"02",x"18",x"1C",x"3A",x"30",x"E1",x"B7", -- 0x25F0
		x"0E",x"D3",x"28",x"0C",x"CB",x"67",x"28",x"06", -- 0x25F8
		x"3A",x"36",x"E1",x"B7",x"20",x"02",x"0E",x"C3", -- 0x2600
		x"3A",x"0E",x"E1",x"B9",x"30",x"BA",x"0E",x"01", -- 0x2608
		x"3A",x"A7",x"E0",x"B1",x"32",x"A7",x"E0",x"3A", -- 0x2610
		x"A7",x"E0",x"B7",x"CA",x"72",x"26",x"08",x"01", -- 0x2618
		x"00",x"01",x"3A",x"99",x"E0",x"FE",x"02",x"30", -- 0x2620
		x"0A",x"08",x"01",x"80",x"01",x"EA",x"33",x"26", -- 0x2628
		x"01",x"00",x"02",x"3A",x"A7",x"E0",x"5F",x"E6", -- 0x2630
		x"03",x"CA",x"54",x"26",x"2A",x"7E",x"E1",x"09", -- 0x2638
		x"54",x"26",x"00",x"22",x"7E",x"E1",x"3A",x"0E", -- 0x2640
		x"E1",x"CB",x"43",x"28",x"03",x"82",x"18",x"01", -- 0x2648
		x"92",x"32",x"0E",x"E1",x"7B",x"E6",x"0C",x"CA", -- 0x2650
		x"72",x"26",x"2A",x"7C",x"E1",x"09",x"54",x"26", -- 0x2658
		x"00",x"22",x"7C",x"E1",x"3A",x"0F",x"E1",x"CB", -- 0x2660
		x"5B",x"28",x"03",x"82",x"18",x"01",x"92",x"32", -- 0x2668
		x"0F",x"E1",x"3A",x"98",x"E0",x"B7",x"20",x"1C", -- 0x2670
		x"3A",x"99",x"E0",x"FE",x"03",x"30",x"15",x"2A", -- 0x2678
		x"0E",x"E1",x"3A",x"97",x"E0",x"FE",x"06",x"38", -- 0x2680
		x"0B",x"FE",x"0B",x"30",x"07",x"7C",x"C6",x"10", -- 0x2688
		x"67",x"22",x"06",x"EB",x"21",x"AE",x"E0",x"3A", -- 0x2690
		x"A7",x"E0",x"4F",x"E6",x"03",x"20",x"15",x"0E", -- 0x2698
		x"03",x"7E",x"E6",x"70",x"FE",x"20",x"3E",x"28", -- 0x26A0
		x"28",x"07",x"34",x"38",x"18",x"35",x"35",x"18", -- 0x26A8
		x"14",x"77",x"18",x"11",x"79",x"E6",x"02",x"7E", -- 0x26B0
		x"20",x"07",x"FE",x"50",x"30",x"07",x"34",x"18", -- 0x26B8
		x"04",x"B7",x"28",x"01",x"35",x"7E",x"B7",x"28", -- 0x26C0
		x"07",x"0F",x"0F",x"0F",x"0F",x"E6",x"07",x"3C", -- 0x26C8
		x"4F",x"06",x"00",x"3A",x"93",x"E0",x"B7",x"20", -- 0x26D0
		x"08",x"21",x"09",x"27",x"09",x"7E",x"32",x"0C", -- 0x26D8
		x"E1",x"3A",x"99",x"E0",x"B7",x"C2",x"3A",x"29", -- 0x26E0
		x"DD",x"21",x"20",x"E1",x"CD",x"F9",x"26",x"DD", -- 0x26E8
		x"21",x"30",x"E1",x"CD",x"F9",x"26",x"C3",x"3A", -- 0x26F0
		x"29",x"DD",x"7E",x"00",x"2F",x"E6",x"82",x"C0", -- 0x26F8
		x"21",x"10",x"27",x"09",x"7E",x"DD",x"77",x"0C", -- 0x2700
		x"C9",x"8C",x"88",x"84",x"80",x"82",x"86",x"8A", -- 0x2708
		x"07",x"24",x"43",x"00",x"34",x"2B",x"01",x"DD", -- 0x2710
		x"21",x"20",x"E1",x"CD",x"22",x"27",x"DD",x"21", -- 0x2718
		x"30",x"E1",x"DD",x"7E",x"00",x"B7",x"C8",x"CB", -- 0x2720
		x"4F",x"CA",x"6A",x"27",x"CB",x"5F",x"C2",x"85", -- 0x2728
		x"28",x"CB",x"57",x"C2",x"6F",x"28",x"2A",x"0E", -- 0x2730
		x"E1",x"CB",x"77",x"3E",x"F3",x"28",x"02",x"3E", -- 0x2738
		x"1D",x"85",x"DD",x"77",x"0E",x"DD",x"7E",x"00", -- 0x2740
		x"E6",x"30",x"20",x"09",x"3A",x"93",x"E0",x"B7", -- 0x2748
		x"20",x"03",x"DD",x"74",x"0F",x"DD",x"35",x"05", -- 0x2750
		x"C2",x"E8",x"2A",x"DD",x"36",x"05",x"02",x"DD", -- 0x2758
		x"7E",x"0D",x"EE",x"01",x"DD",x"77",x"0D",x"C3", -- 0x2760
		x"E8",x"2A",x"CB",x"7F",x"C8",x"DD",x"7E",x"01", -- 0x2768
		x"CD",x"F7",x"66",x"7D",x"27",x"99",x"27",x"D4", -- 0x2770
		x"27",x"08",x"28",x"1D",x"28",x"CD",x"D6",x"28", -- 0x2778
		x"DD",x"36",x"0D",x"12",x"DD",x"36",x"0F",x"00", -- 0x2780
		x"DD",x"36",x"0C",x"20",x"DD",x"36",x"05",x"02", -- 0x2788
		x"DD",x"36",x"07",x"08",x"DD",x"34",x"01",x"18", -- 0x2790
		x"BC",x"CD",x"D6",x"28",x"01",x"FC",x"FF",x"3A", -- 0x2798
		x"0F",x"E1",x"C6",x"18",x"DD",x"BE",x"0F",x"38", -- 0x27A0
		x"03",x"01",x"FE",x"FF",x"CD",x"09",x"62",x"09", -- 0x27A8
		x"CD",x"C8",x"50",x"CD",x"5A",x"28",x"DD",x"CB", -- 0x27B0
		x"0D",x"66",x"20",x"99",x"3A",x"0F",x"E1",x"C6", -- 0x27B8
		x"10",x"4F",x"DD",x"7E",x"0F",x"91",x"30",x"8D", -- 0x27C0
		x"AF",x"DD",x"77",x"02",x"CD",x"3C",x"28",x"DD", -- 0x27C8
		x"34",x"01",x"18",x"81",x"CD",x"5A",x"28",x"DD", -- 0x27D0
		x"35",x"03",x"20",x"12",x"DD",x"34",x"02",x"CD", -- 0x27D8
		x"3C",x"28",x"30",x"0A",x"DD",x"34",x"01",x"DD", -- 0x27E0
		x"36",x"02",x"00",x"CD",x"41",x"28",x"DD",x"4E", -- 0x27E8
		x"04",x"CB",x"79",x"06",x"00",x"28",x"01",x"05", -- 0x27F0
		x"3A",x"0F",x"E1",x"6F",x"26",x"00",x"09",x"CD", -- 0x27F8
		x"C8",x"50",x"CD",x"D6",x"28",x"C3",x"55",x"27", -- 0x2800
		x"CD",x"5A",x"28",x"DD",x"35",x"03",x"20",x"DE", -- 0x2808
		x"DD",x"34",x"02",x"CD",x"41",x"28",x"30",x"D6", -- 0x2810
		x"DD",x"34",x"01",x"18",x"D1",x"CD",x"5A",x"28", -- 0x2818
		x"CD",x"D6",x"28",x"3A",x"0F",x"E1",x"DD",x"77", -- 0x2820
		x"0F",x"DD",x"7E",x"07",x"B7",x"C2",x"EE",x"27", -- 0x2828
		x"DD",x"7E",x"00",x"E6",x"F3",x"F6",x"02",x"DD", -- 0x2830
		x"77",x"00",x"18",x"B2",x"21",x"4C",x"87",x"18", -- 0x2838
		x"03",x"21",x"53",x"87",x"DD",x"7E",x"02",x"07", -- 0x2840
		x"4F",x"06",x"00",x"09",x"7E",x"B7",x"3F",x"C8", -- 0x2848
		x"DD",x"77",x"03",x"23",x"7E",x"DD",x"77",x"04", -- 0x2850
		x"B7",x"C9",x"DD",x"7E",x"07",x"3C",x"E6",x"0F", -- 0x2858
		x"DD",x"77",x"07",x"21",x"D4",x"78",x"4F",x"06", -- 0x2860
		x"00",x"09",x"7E",x"DD",x"77",x"0C",x"C9",x"AF", -- 0x2868
		x"DD",x"77",x"02",x"DD",x"CB",x"00",x"DE",x"DD", -- 0x2870
		x"36",x"0C",x"D8",x"DD",x"36",x"0D",x"0E",x"CD", -- 0x2878
		x"BD",x"28",x"C3",x"E8",x"2A",x"DD",x"35",x"03", -- 0x2880
		x"C0",x"DD",x"34",x"02",x"CD",x"BD",x"28",x"D2", -- 0x2888
		x"E8",x"2A",x"DD",x"36",x"0D",x"10",x"DD",x"77", -- 0x2890
		x"0E",x"DD",x"77",x"0F",x"CD",x"E8",x"2A",x"DD", -- 0x2898
		x"7E",x"0B",x"CD",x"05",x"67",x"DD",x"36",x"00", -- 0x28A0
		x"00",x"3A",x"20",x"E1",x"4F",x"3A",x"30",x"E1", -- 0x28A8
		x"B1",x"E6",x"80",x"C0",x"3A",x"1F",x"E1",x"E6", -- 0x28B0
		x"FE",x"32",x"1F",x"E1",x"C9",x"DD",x"7E",x"02", -- 0x28B8
		x"07",x"4F",x"06",x"00",x"21",x"87",x"87",x"09", -- 0x28C0
		x"7E",x"B7",x"37",x"C8",x"DD",x"77",x"03",x"23", -- 0x28C8
		x"7E",x"DD",x"77",x"0C",x"B7",x"C9",x"DD",x"CB", -- 0x28D0
		x"00",x"76",x"3A",x"0E",x"E1",x"06",x"F3",x"28", -- 0x28D8
		x"02",x"06",x"1D",x"80",x"DD",x"77",x"0E",x"C9", -- 0x28E0
		x"3A",x"20",x"E1",x"0F",x"38",x"0E",x"DD",x"21", -- 0x28E8
		x"20",x"E1",x"CD",x"23",x"29",x"38",x"05",x"21", -- 0x28F0
		x"18",x"E1",x"CB",x"86",x"3A",x"30",x"E1",x"0F", -- 0x28F8
		x"38",x"0E",x"DD",x"21",x"30",x"E1",x"CD",x"23", -- 0x2900
		x"29",x"38",x"05",x"21",x"18",x"E1",x"CB",x"8E", -- 0x2908
		x"3A",x"18",x"E1",x"E6",x"03",x"C0",x"21",x"20", -- 0x2910
		x"E1",x"CB",x"FE",x"21",x"30",x"E1",x"CB",x"FE", -- 0x2918
		x"CB",x"F6",x"C9",x"16",x"03",x"CD",x"51",x"0C", -- 0x2920
		x"D8",x"7D",x"E6",x"1F",x"07",x"07",x"DD",x"77", -- 0x2928
		x"0B",x"DD",x"36",x"00",x"01",x"AF",x"DD",x"77", -- 0x2930
		x"01",x"C9",x"21",x"0C",x"E1",x"11",x"00",x"EB", -- 0x2938
		x"01",x"04",x"00",x"ED",x"B0",x"C9",x"06",x"03", -- 0x2940
		x"DD",x"21",x"60",x"E2",x"11",x"10",x"00",x"21", -- 0x2948
		x"A1",x"E0",x"DD",x"CB",x"00",x"46",x"28",x"05", -- 0x2950
		x"DD",x"19",x"10",x"F6",x"C9",x"34",x"2A",x"0E", -- 0x2958
		x"E1",x"06",x"BC",x"0E",x"4E",x"3A",x"64",x"E1", -- 0x2960
		x"07",x"7D",x"38",x"06",x"C6",x"08",x"06",x"BA", -- 0x2968
		x"0E",x"0E",x"DD",x"77",x"0E",x"7C",x"C6",x"0B", -- 0x2970
		x"DD",x"77",x"0F",x"DD",x"70",x"0C",x"DD",x"71", -- 0x2978
		x"0D",x"0E",x"00",x"3A",x"30",x"E1",x"CB",x"67", -- 0x2980
		x"20",x"08",x"E6",x"8E",x"FE",x"82",x"20",x"02", -- 0x2988
		x"0E",x"10",x"3A",x"20",x"E1",x"CB",x"67",x"20", -- 0x2990
		x"08",x"E6",x"8E",x"FE",x"82",x"20",x"02",x"CB", -- 0x2998
		x"E9",x"DD",x"36",x"01",x"00",x"DD",x"7E",x"00", -- 0x29A0
		x"E6",x"80",x"3C",x"B1",x"DD",x"77",x"00",x"79", -- 0x29A8
		x"B7",x"C8",x"FD",x"21",x"20",x"E1",x"CD",x"BD", -- 0x29B0
		x"29",x"FD",x"21",x"30",x"E1",x"FD",x"7E",x"00", -- 0x29B8
		x"4F",x"2F",x"E6",x"82",x"C0",x"79",x"E6",x"0C", -- 0x29C0
		x"C0",x"79",x"CB",x"77",x"01",x"30",x"00",x"28", -- 0x29C8
		x"03",x"01",x"60",x"00",x"DD",x"E5",x"DD",x"09", -- 0x29D0
		x"4F",x"06",x"01",x"FD",x"7E",x"0E",x"5F",x"FE", -- 0x29D8
		x"7A",x"30",x"0E",x"04",x"FE",x"77",x"38",x"09", -- 0x29E0
		x"1E",x"76",x"CB",x"71",x"28",x"03",x"1E",x"7A", -- 0x29E8
		x"05",x"DD",x"56",x"04",x"CB",x"40",x"28",x"03", -- 0x29F0
		x"DD",x"56",x"05",x"DD",x"72",x"0B",x"DD",x"36", -- 0x29F8
		x"0C",x"B9",x"DD",x"36",x"0D",x"0E",x"DD",x"73", -- 0x2A00
		x"0E",x"FD",x"7E",x"0F",x"C6",x"0B",x"DD",x"77", -- 0x2A08
		x"0F",x"79",x"E6",x"40",x"F6",x"81",x"DD",x"77", -- 0x2A10
		x"00",x"DD",x"E1",x"C9",x"DD",x"CB",x"01",x"46", -- 0x2A18
		x"C2",x"43",x"2A",x"CB",x"5F",x"C2",x"9C",x"2A", -- 0x2A20
		x"CB",x"57",x"C2",x"6A",x"2A",x"DD",x"7E",x"0F", -- 0x2A28
		x"C6",x"06",x"38",x"0F",x"DD",x"77",x"0F",x"DD", -- 0x2A30
		x"77",x"3F",x"DD",x"77",x"6F",x"CD",x"C5",x"2A", -- 0x2A38
		x"C3",x"AC",x"1C",x"AF",x"DD",x"77",x"0D",x"DD", -- 0x2A40
		x"77",x"0E",x"DD",x"7E",x"00",x"E6",x"30",x"28", -- 0x2A48
		x"0C",x"CD",x"F9",x"2A",x"CD",x"C5",x"2A",x"AF", -- 0x2A50
		x"DD",x"77",x"00",x"18",x"07",x"DD",x"36",x"00", -- 0x2A58
		x"00",x"CD",x"E8",x"2A",x"CD",x"BD",x"2A",x"C3", -- 0x2A60
		x"AC",x"1C",x"DD",x"CB",x"0D",x"76",x"CA",x"79", -- 0x2A68
		x"2A",x"DD",x"7E",x"0E",x"C6",x"08",x"DD",x"77", -- 0x2A70
		x"0E",x"DD",x"36",x"0C",x"D8",x"DD",x"36",x"0D", -- 0x2A78
		x"0E",x"DD",x"36",x"0A",x"00",x"DD",x"CB",x"00", -- 0x2A80
		x"DE",x"DD",x"7E",x"00",x"E6",x"30",x"C4",x"F9", -- 0x2A88
		x"2A",x"CD",x"C5",x"2A",x"0E",x"03",x"CD",x"78", -- 0x2A90
		x"11",x"C3",x"AC",x"1C",x"DD",x"34",x"0A",x"DD", -- 0x2A98
		x"7E",x"0A",x"FE",x"06",x"D2",x"AD",x"2A",x"DD", -- 0x2AA0
		x"34",x"0C",x"C3",x"B7",x"2A",x"AF",x"DD",x"77", -- 0x2AA8
		x"0E",x"DD",x"77",x"00",x"CD",x"BD",x"2A",x"CD", -- 0x2AB0
		x"E8",x"2A",x"C3",x"AC",x"1C",x"21",x"A1",x"E0", -- 0x2AB8
		x"7E",x"B7",x"C8",x"35",x"C9",x"DD",x"4E",x"00", -- 0x2AC0
		x"79",x"E6",x"30",x"CA",x"E8",x"2A",x"DD",x"E5", -- 0x2AC8
		x"E1",x"C5",x"01",x"3B",x"00",x"09",x"CB",x"6F", -- 0x2AD0
		x"C4",x"EF",x"2A",x"C1",x"DD",x"E5",x"E1",x"CB", -- 0x2AD8
		x"61",x"01",x"6B",x"00",x"09",x"C4",x"EF",x"2A", -- 0x2AE0
		x"DD",x"E5",x"E1",x"01",x"0B",x"00",x"09",x"5E", -- 0x2AE8
		x"23",x"16",x"EB",x"01",x"04",x"00",x"ED",x"B0", -- 0x2AF0
		x"C9",x"AF",x"DD",x"77",x"30",x"DD",x"77",x"3E", -- 0x2AF8
		x"DD",x"77",x"60",x"DD",x"77",x"6E",x"C9",x"AF", -- 0x2B00
		x"32",x"41",x"E1",x"21",x"B4",x"A8",x"22",x"58", -- 0x2B08
		x"E1",x"CD",x"44",x"2B",x"CD",x"68",x"2B",x"06", -- 0x2B10
		x"0A",x"C5",x"06",x"01",x"DF",x"3A",x"A4",x"E9", -- 0x2B18
		x"B7",x"C4",x"8A",x"2B",x"C1",x"10",x"F2",x"3A", -- 0x2B20
		x"41",x"E1",x"3C",x"FE",x"06",x"38",x"01",x"AF", -- 0x2B28
		x"32",x"41",x"E1",x"20",x"DF",x"3A",x"40",x"E1", -- 0x2B30
		x"3C",x"FE",x"80",x"38",x"02",x"3E",x"40",x"32", -- 0x2B38
		x"40",x"E1",x"18",x"C7",x"3A",x"40",x"E1",x"6F", -- 0x2B40
		x"26",x"00",x"29",x"29",x"EB",x"2A",x"58",x"E1", -- 0x2B48
		x"19",x"7E",x"32",x"52",x"E1",x"23",x"7E",x"32", -- 0x2B50
		x"51",x"E1",x"E6",x"80",x"32",x"43",x"E1",x"23", -- 0x2B58
		x"4E",x"23",x"46",x"ED",x"43",x"72",x"E1",x"C9", -- 0x2B60
		x"3A",x"51",x"E1",x"CB",x"7F",x"28",x"09",x"CB", -- 0x2B68
		x"77",x"20",x"13",x"3A",x"52",x"E1",x"18",x"0A", -- 0x2B70
		x"57",x"3A",x"52",x"E1",x"5F",x"3A",x"E8",x"E0", -- 0x2B78
		x"A3",x"82",x"32",x"53",x"E1",x"AF",x"32",x"43", -- 0x2B80
		x"E1",x"C9",x"DD",x"2A",x"A0",x"E9",x"FD",x"21", -- 0x2B88
		x"00",x"E7",x"AF",x"F3",x"FD",x"36",x"00",x"FF", -- 0x2B90
		x"32",x"45",x"E1",x"FB",x"21",x"06",x"C8",x"F3", -- 0x2B98
		x"36",x"01",x"DD",x"56",x"00",x"DD",x"46",x"01", -- 0x2BA0
		x"36",x"00",x"FB",x"7A",x"FE",x"FF",x"CA",x"BF", -- 0x2BA8
		x"2C",x"FE",x"FD",x"28",x"1B",x"FE",x"FC",x"20", -- 0x2BB0
		x"05",x"32",x"C7",x"E0",x"18",x"12",x"FE",x"FE", -- 0x2BB8
		x"CA",x"BD",x"2C",x"CB",x"7F",x"28",x"37",x"CB", -- 0x2BC0
		x"77",x"20",x"09",x"E6",x"0F",x"32",x"71",x"E1", -- 0x2BC8
		x"DD",x"23",x"18",x"C8",x"4F",x"E6",x"0F",x"57", -- 0x2BD0
		x"3A",x"04",x"C0",x"CB",x"77",x"7A",x"20",x"02", -- 0x2BD8
		x"C6",x"02",x"32",x"6B",x"E1",x"79",x"0F",x"0F", -- 0x2BE0
		x"0F",x"0F",x"E6",x"03",x"4F",x"28",x"07",x"3A", -- 0x2BE8
		x"C5",x"E0",x"B7",x"28",x"01",x"0D",x"79",x"32", -- 0x2BF0
		x"6A",x"E1",x"DD",x"23",x"18",x"9E",x"7A",x"E6", -- 0x2BF8
		x"1F",x"FE",x"08",x"20",x"1C",x"3A",x"05",x"EC", -- 0x2C00
		x"B7",x"C2",x"B3",x"2C",x"7A",x"07",x"07",x"07", -- 0x2C08
		x"E6",x"03",x"F6",x"80",x"32",x"00",x"EC",x"32", -- 0x2C10
		x"05",x"EC",x"78",x"32",x"22",x"EC",x"C3",x"B3", -- 0x2C18
		x"2C",x"FE",x"09",x"20",x"16",x"78",x"E6",x"01", -- 0x2C20
		x"07",x"07",x"07",x"4F",x"7A",x"07",x"07",x"07", -- 0x2C28
		x"E6",x"03",x"F6",x"80",x"B1",x"32",x"B0",x"E7", -- 0x2C30
		x"C3",x"B3",x"2C",x"FE",x"10",x"20",x"1E",x"3A", -- 0x2C38
		x"E0",x"E7",x"B7",x"20",x"6E",x"78",x"E6",x"0F", -- 0x2C40
		x"FE",x"04",x"20",x"08",x"3A",x"13",x"E1",x"B7", -- 0x2C48
		x"3E",x"04",x"20",x"5F",x"F6",x"80",x"6F",x"60", -- 0x2C50
		x"22",x"E0",x"E7",x"18",x"56",x"FE",x"03",x"28", -- 0x2C58
		x"43",x"FE",x"04",x"28",x"12",x"FD",x"70",x"01", -- 0x2C60
		x"FD",x"36",x"02",x"FF",x"21",x"45",x"E1",x"F3", -- 0x2C68
		x"FD",x"72",x"00",x"34",x"FB",x"18",x"3C",x"CB", -- 0x2C70
		x"70",x"78",x"20",x"22",x"E6",x"30",x"0F",x"0F", -- 0x2C78
		x"0F",x"0F",x"32",x"1C",x"E1",x"78",x"E6",x"0F", -- 0x2C80
		x"47",x"21",x"1B",x"E1",x"F3",x"32",x"1D",x"E1", -- 0x2C88
		x"3A",x"1E",x"E1",x"B7",x"20",x"05",x"78",x"77", -- 0x2C90
		x"32",x"1E",x"E1",x"FB",x"18",x"15",x"AF",x"32", -- 0x2C98
		x"1D",x"E1",x"18",x"0F",x"3A",x"14",x"E1",x"B7", -- 0x2CA0
		x"20",x"09",x"7A",x"E6",x"60",x"3C",x"4F",x"ED", -- 0x2CA8
		x"43",x"14",x"E1",x"01",x"02",x"00",x"FD",x"09", -- 0x2CB0
		x"DD",x"09",x"C3",x"9C",x"2B",x"DD",x"23",x"DD", -- 0x2CB8
		x"22",x"A0",x"E9",x"FD",x"36",x"00",x"FF",x"AF", -- 0x2CC0
		x"32",x"A4",x"E9",x"C9",x"DD",x"7E",x"00",x"B7", -- 0x2CC8
		x"C8",x"4F",x"DD",x"46",x"01",x"DD",x"6E",x"02", -- 0x2CD0
		x"DD",x"66",x"03",x"DD",x"56",x"04",x"CD",x"53", -- 0x2CD8
		x"02",x"0E",x"05",x"DD",x"09",x"18",x"E5",x"06", -- 0x2CE0
		x"05",x"3E",x"01",x"EF",x"3C",x"10",x"FC",x"3E", -- 0x2CE8
		x"07",x"EF",x"3C",x"EF",x"3C",x"EF",x"3E",x"0B", -- 0x2CF0
		x"EF",x"3E",x"0D",x"EF",x"C9",x"21",x"D4",x"E0", -- 0x2CF8
		x"CB",x"E6",x"7E",x"32",x"04",x"C8",x"CB",x"A6", -- 0x2D00
		x"F3",x"3A",x"D4",x"E0",x"32",x"04",x"C8",x"FB", -- 0x2D08
		x"C9",x"06",x"08",x"AF",x"77",x"23",x"10",x"FC", -- 0x2D10
		x"C9",x"DD",x"56",x"00",x"DD",x"4E",x"01",x"DD", -- 0x2D18
		x"46",x"02",x"DD",x"7E",x"03",x"FF",x"01",x"03", -- 0x2D20
		x"00",x"DD",x"09",x"15",x"20",x"EE",x"C9",x"3A", -- 0x2D28
		x"A6",x"E0",x"E6",x"02",x"C9",x"3A",x"00",x"E0", -- 0x2D30
		x"07",x"D2",x"41",x"11",x"3A",x"03",x"C0",x"E6", -- 0x2D38
		x"08",x"3A",x"01",x"C0",x"28",x"0B",x"CD",x"2F", -- 0x2D40
		x"2D",x"3A",x"01",x"C0",x"28",x"03",x"3A",x"02", -- 0x2D48
		x"C0",x"2F",x"E6",x"3F",x"C9",x"3A",x"00",x"E0", -- 0x2D50
		x"07",x"D0",x"ED",x"5B",x"4A",x"E0",x"ED",x"4B", -- 0x2D58
		x"48",x"E0",x"CD",x"2F",x"2D",x"28",x"08",x"ED", -- 0x2D60
		x"5B",x"52",x"E0",x"ED",x"4B",x"50",x"E0",x"79", -- 0x2D68
		x"B7",x"C2",x"D3",x"2D",x"B0",x"C0",x"2A",x"10", -- 0x2D70
		x"E1",x"7B",x"BD",x"38",x"2A",x"20",x"04",x"7A", -- 0x2D78
		x"BC",x"38",x"24",x"3A",x"03",x"C0",x"E6",x"10", -- 0x2D80
		x"11",x"00",x"08",x"20",x"03",x"11",x"01",x"00", -- 0x2D88
		x"7A",x"84",x"FE",x"0A",x"38",x"03",x"D6",x"0A", -- 0x2D90
		x"2C",x"67",x"7B",x"85",x"6F",x"22",x"10",x"E1", -- 0x2D98
		x"21",x"01",x"E1",x"34",x"CD",x"C9",x"2D",x"3A", -- 0x2DA0
		x"00",x"E1",x"E6",x"02",x"C0",x"7A",x"53",x"5F", -- 0x2DA8
		x"3A",x"03",x"C0",x"E6",x"20",x"21",x"FE",x"FF", -- 0x2DB0
		x"20",x"01",x"2D",x"19",x"D0",x"3A",x"00",x"E1", -- 0x2DB8
		x"F6",x"02",x"32",x"00",x"E1",x"21",x"01",x"E1", -- 0x2DC0
		x"34",x"0E",x"08",x"CD",x"78",x"11",x"CD",x"6D", -- 0x2DC8
		x"12",x"AF",x"C9",x"21",x"48",x"E0",x"CD",x"2F", -- 0x2DD0
		x"2D",x"0E",x"0A",x"28",x"05",x"0E",x"0F",x"21", -- 0x2DD8
		x"50",x"E0",x"3E",x"01",x"77",x"23",x"06",x"07", -- 0x2DE0
		x"CD",x"13",x"2D",x"CD",x"14",x"13",x"AF",x"01", -- 0x2DE8
		x"F7",x"6F",x"FF",x"37",x"C9",x"DD",x"21",x"00", -- 0x2DF0
		x"E4",x"06",x"10",x"DD",x"CB",x"00",x"46",x"C2", -- 0x2DF8
		x"F3",x"2E",x"11",x"30",x"00",x"DD",x"19",x"10", -- 0x2E00
		x"F2",x"DD",x"21",x"00",x"E3",x"3A",x"F0",x"E3", -- 0x2E08
		x"47",x"0E",x"0F",x"C5",x"DD",x"7E",x"00",x"CB", -- 0x2E10
		x"47",x"CA",x"B0",x"2E",x"CB",x"67",x"C2",x"DF", -- 0x2E18
		x"2E",x"CB",x"5F",x"C2",x"C4",x"2E",x"CB",x"4F", -- 0x2E20
		x"C2",x"B0",x"2E",x"C1",x"05",x"C5",x"CB",x"57", -- 0x2E28
		x"C2",x"A5",x"2E",x"DD",x"56",x"09",x"DD",x"4E", -- 0x2E30
		x"05",x"DD",x"46",x"06",x"DD",x"6E",x"03",x"26", -- 0x2E38
		x"00",x"09",x"DD",x"75",x"03",x"DD",x"7E",x"0E", -- 0x2E40
		x"CB",x"42",x"20",x"03",x"84",x"18",x"01",x"94", -- 0x2E48
		x"DA",x"A5",x"2E",x"DD",x"77",x"0E",x"DD",x"4E", -- 0x2E50
		x"07",x"DD",x"46",x"08",x"DD",x"6E",x"04",x"26", -- 0x2E58
		x"00",x"09",x"DD",x"75",x"04",x"DD",x"7E",x"0F", -- 0x2E60
		x"CB",x"4A",x"20",x"03",x"84",x"18",x"01",x"94", -- 0x2E68
		x"DD",x"77",x"0F",x"D2",x"7A",x"2E",x"DD",x"CB", -- 0x2E70
		x"0D",x"E6",x"DD",x"CB",x"0D",x"66",x"CA",x"86", -- 0x2E78
		x"2E",x"FE",x"F0",x"DA",x"A5",x"2E",x"CD",x"E8", -- 0x2E80
		x"2A",x"CD",x"B6",x"38",x"30",x"17",x"3A",x"A5", -- 0x2E88
		x"E0",x"B7",x"20",x"1C",x"CD",x"94",x"38",x"38", -- 0x2E90
		x"17",x"3E",x"01",x"32",x"A5",x"E0",x"AF",x"01", -- 0x2E98
		x"30",x"67",x"FF",x"18",x"00",x"21",x"F0",x"E3", -- 0x2EA0
		x"35",x"CD",x"94",x"61",x"DD",x"36",x"00",x"00", -- 0x2EA8
		x"01",x"10",x"00",x"DD",x"09",x"C1",x"78",x"B7", -- 0x2EB0
		x"28",x"04",x"0D",x"C2",x"13",x"2E",x"06",x"01", -- 0x2EB8
		x"DF",x"C3",x"F5",x"2D",x"DD",x"36",x"0C",x"D8", -- 0x2EC0
		x"DD",x"36",x"0D",x"0E",x"DD",x"36",x"0A",x"00", -- 0x2EC8
		x"DD",x"CB",x"00",x"E6",x"CD",x"E8",x"2A",x"0E", -- 0x2ED0
		x"03",x"CD",x"78",x"11",x"C3",x"B0",x"2E",x"DD", -- 0x2ED8
		x"34",x"0A",x"DD",x"7E",x"0A",x"FE",x"06",x"D2", -- 0x2EE0
		x"A5",x"2E",x"DD",x"34",x"0C",x"CD",x"E8",x"2A", -- 0x2EE8
		x"C3",x"B0",x"2E",x"C5",x"DD",x"7E",x"00",x"CB", -- 0x2EF0
		x"4F",x"C2",x"27",x"62",x"07",x"07",x"E6",x"03", -- 0x2EF8
		x"CA",x"27",x"2F",x"3D",x"CA",x"14",x"30",x"3D", -- 0x2F00
		x"CA",x"E4",x"30",x"11",x"47",x"2F",x"D5",x"DD", -- 0x2F08
		x"7E",x"03",x"E6",x"07",x"CD",x"F7",x"66",x"FE", -- 0x2F10
		x"51",x"40",x"52",x"67",x"52",x"67",x"52",x"B8", -- 0x2F18
		x"52",x"F2",x"52",x"C1",x"C3",x"02",x"2E",x"DD", -- 0x2F20
		x"7E",x"01",x"07",x"07",x"E6",x"03",x"C2",x"5D", -- 0x2F28
		x"2F",x"11",x"47",x"2F",x"D5",x"DD",x"7E",x"03", -- 0x2F30
		x"E6",x"03",x"CA",x"F3",x"30",x"3D",x"CA",x"51", -- 0x2F38
		x"31",x"CD",x"25",x"33",x"C3",x"54",x"32",x"DD", -- 0x2F40
		x"7E",x"18",x"EE",x"01",x"DD",x"77",x"18",x"E6", -- 0x2F48
		x"01",x"20",x"D0",x"DD",x"7E",x"0D",x"EE",x"01", -- 0x2F50
		x"DD",x"77",x"0D",x"18",x"C6",x"3D",x"C2",x"8C", -- 0x2F58
		x"2F",x"11",x"23",x"2F",x"D5",x"DD",x"7E",x"03", -- 0x2F60
		x"E6",x"03",x"CA",x"7A",x"2F",x"3D",x"CA",x"59", -- 0x2F68
		x"31",x"CD",x"25",x"33",x"CD",x"25",x"34",x"C3", -- 0x2F70
		x"2A",x"4B",x"CD",x"82",x"36",x"DD",x"36",x"0A", -- 0x2F78
		x"00",x"CD",x"37",x"31",x"D6",x"03",x"CA",x"C6", -- 0x2F80
		x"3E",x"C3",x"E6",x"3E",x"3D",x"C2",x"BA",x"2F", -- 0x2F88
		x"CD",x"25",x"33",x"11",x"23",x"2F",x"D5",x"DD", -- 0x2F90
		x"7E",x"03",x"E6",x"0F",x"F5",x"C4",x"25",x"34", -- 0x2F98
		x"F1",x"CD",x"F7",x"66",x"49",x"47",x"EE",x"47", -- 0x2FA0
		x"4E",x"48",x"63",x"48",x"91",x"48",x"03",x"49", -- 0x2FA8
		x"9B",x"49",x"BD",x"49",x"00",x"4A",x"48",x"4A", -- 0x2FB0
		x"7D",x"4A",x"11",x"CF",x"2F",x"D5",x"CD",x"7E", -- 0x2FB8
		x"33",x"DD",x"7E",x"03",x"E6",x"03",x"CA",x"6A", -- 0x2FC0
		x"4E",x"CD",x"25",x"34",x"C3",x"26",x"4F",x"DD", -- 0x2FC8
		x"7E",x"18",x"EE",x"01",x"DD",x"77",x"18",x"E6", -- 0x2FD0
		x"01",x"C2",x"EC",x"2F",x"DD",x"7E",x"0D",x"EE", -- 0x2FD8
		x"01",x"DD",x"77",x"0D",x"DD",x"7E",x"2D",x"EE", -- 0x2FE0
		x"01",x"DD",x"77",x"2D",x"DD",x"7E",x"18",x"CB", -- 0x2FE8
		x"4F",x"CA",x"23",x"2F",x"C6",x"20",x"DD",x"77", -- 0x2FF0
		x"18",x"D2",x"23",x"2F",x"F6",x"20",x"DD",x"77", -- 0x2FF8
		x"18",x"16",x"02",x"DD",x"7E",x"0D",x"AA",x"DD", -- 0x3000
		x"77",x"0D",x"DD",x"7E",x"2D",x"AA",x"DD",x"77", -- 0x3008
		x"2D",x"C3",x"23",x"2F",x"DD",x"CB",x"01",x"76", -- 0x3010
		x"C2",x"80",x"30",x"11",x"34",x"30",x"D5",x"DD", -- 0x3018
		x"7E",x"03",x"E6",x"03",x"CA",x"F9",x"52",x"3D", -- 0x3020
		x"CA",x"30",x"54",x"CD",x"4C",x"33",x"CD",x"25", -- 0x3028
		x"34",x"C3",x"51",x"54",x"DD",x"7E",x"18",x"EE", -- 0x3030
		x"01",x"DD",x"77",x"18",x"E6",x"01",x"C2",x"4A", -- 0x3038
		x"30",x"16",x"01",x"3A",x"18",x"EC",x"AA",x"32", -- 0x3040
		x"18",x"EC",x"DD",x"7E",x"18",x"CB",x"4F",x"CA", -- 0x3048
		x"23",x"2F",x"C6",x"20",x"DD",x"77",x"18",x"D2", -- 0x3050
		x"23",x"2F",x"F6",x"20",x"DD",x"77",x"18",x"16", -- 0x3058
		x"02",x"DD",x"7E",x"0D",x"AA",x"DD",x"77",x"0D", -- 0x3060
		x"3A",x"13",x"EC",x"AA",x"32",x"13",x"EC",x"3A", -- 0x3068
		x"18",x"EC",x"AA",x"32",x"18",x"EC",x"3A",x"1D", -- 0x3070
		x"EC",x"AA",x"32",x"1D",x"EC",x"C3",x"23",x"2F", -- 0x3078
		x"11",x"99",x"30",x"D5",x"DD",x"7E",x"03",x"E6", -- 0x3080
		x"03",x"CA",x"31",x"59",x"3D",x"C2",x"3C",x"5A", -- 0x3088
		x"CD",x"BA",x"30",x"CD",x"25",x"34",x"C3",x"F4", -- 0x3090
		x"59",x"DD",x"7E",x"18",x"EE",x"80",x"DD",x"77", -- 0x3098
		x"18",x"4F",x"E6",x"80",x"C2",x"23",x"2F",x"16", -- 0x30A0
		x"01",x"3A",x"59",x"EB",x"AA",x"32",x"59",x"EB", -- 0x30A8
		x"3A",x"79",x"EB",x"AA",x"32",x"79",x"EB",x"C3", -- 0x30B0
		x"23",x"2F",x"3A",x"99",x"E0",x"B7",x"C0",x"21", -- 0x30B8
		x"D4",x"37",x"DD",x"E5",x"FD",x"E1",x"CD",x"6C", -- 0x30C0
		x"37",x"30",x"05",x"CD",x"96",x"33",x"30",x"0F", -- 0x30C8
		x"21",x"D8",x"37",x"DD",x"E5",x"FD",x"E1",x"CD", -- 0x30D0
		x"A0",x"37",x"D0",x"CD",x"96",x"33",x"D8",x"B7", -- 0x30D8
		x"CA",x"41",x"33",x"C9",x"11",x"23",x"2F",x"D5", -- 0x30E0
		x"DD",x"7E",x"03",x"E6",x"03",x"CA",x"BA",x"5F", -- 0x30E8
		x"C3",x"A1",x"61",x"CD",x"82",x"36",x"DD",x"36", -- 0x30F0
		x"18",x"01",x"DD",x"36",x"0A",x"00",x"DD",x"7E", -- 0x30F8
		x"08",x"E6",x"E0",x"20",x"2B",x"DD",x"4E",x"1A", -- 0x3100
		x"06",x"00",x"21",x"34",x"31",x"09",x"DD",x"7E", -- 0x3108
		x"0D",x"E6",x"F0",x"B6",x"DD",x"77",x"0D",x"DD", -- 0x3110
		x"CB",x"01",x"6E",x"C2",x"3B",x"42",x"CD",x"37", -- 0x3118
		x"31",x"CD",x"F7",x"66",x"FA",x"38",x"94",x"3B", -- 0x3120
		x"1B",x"3D",x"30",x"3D",x"2A",x"3E",x"2A",x"41", -- 0x3128
		x"DD",x"34",x"03",x"C9",x"00",x"02",x"04",x"DD", -- 0x3130
		x"7E",x"05",x"07",x"4F",x"06",x"00",x"21",x"80", -- 0x3138
		x"A7",x"09",x"4E",x"23",x"46",x"0A",x"DD",x"77", -- 0x3140
		x"12",x"03",x"DD",x"71",x"10",x"DD",x"70",x"11", -- 0x3148
		x"C9",x"DD",x"7E",x"08",x"E6",x"E0",x"C2",x"97", -- 0x3150
		x"31",x"DD",x"CB",x"01",x"6E",x"C2",x"B3",x"43", -- 0x3158
		x"21",x"7C",x"79",x"DD",x"7E",x"14",x"07",x"4F", -- 0x3160
		x"06",x"00",x"CD",x"E0",x"3C",x"0E",x"02",x"DD", -- 0x3168
		x"7E",x"0D",x"CB",x"67",x"20",x"01",x"0C",x"79", -- 0x3170
		x"FE",x"03",x"C2",x"E8",x"2A",x"01",x"E8",x"2A", -- 0x3178
		x"C5",x"AF",x"DD",x"77",x"13",x"DD",x"7E",x"12", -- 0x3180
		x"CD",x"F7",x"66",x"24",x"39",x"B2",x"3B",x"A9", -- 0x3188
		x"3B",x"06",x"3F",x"2D",x"3F",x"72",x"41",x"E6", -- 0x3190
		x"C0",x"FE",x"80",x"CA",x"30",x"32",x"DD",x"7E", -- 0x3198
		x"14",x"B7",x"28",x"04",x"DD",x"35",x"14",x"C9", -- 0x31A0
		x"CD",x"DE",x"31",x"DD",x"35",x"13",x"20",x"04", -- 0x31A8
		x"DD",x"36",x"03",x"02",x"DD",x"7E",x"0D",x"E6", -- 0x31B0
		x"10",x"C2",x"E8",x"2A",x"DD",x"CB",x"00",x"A6", -- 0x31B8
		x"DD",x"CB",x"02",x"E6",x"DD",x"7E",x"08",x"E6", -- 0x31C0
		x"E0",x"FE",x"60",x"CA",x"E8",x"2A",x"DD",x"7E", -- 0x31C8
		x"02",x"E6",x"0F",x"FE",x"04",x"C2",x"E8",x"2A", -- 0x31D0
		x"32",x"13",x"E1",x"C3",x"E8",x"2A",x"DD",x"6E", -- 0x31D8
		x"10",x"DD",x"66",x"11",x"4E",x"23",x"7E",x"DD", -- 0x31E0
		x"CB",x"02",x"6E",x"28",x"02",x"ED",x"44",x"47", -- 0x31E8
		x"C3",x"E4",x"3C",x"DD",x"6E",x"10",x"DD",x"66", -- 0x31F0
		x"11",x"DD",x"7E",x"0F",x"86",x"DD",x"77",x"0F", -- 0x31F8
		x"CB",x"7E",x"20",x"01",x"3F",x"DD",x"7E",x"0D", -- 0x3200
		x"38",x"05",x"EE",x"10",x"DD",x"77",x"0D",x"CB", -- 0x3208
		x"67",x"28",x"06",x"DD",x"7E",x"0F",x"FE",x"F1", -- 0x3210
		x"D8",x"23",x"7E",x"DD",x"CB",x"02",x"6E",x"28", -- 0x3218
		x"02",x"ED",x"44",x"47",x"DD",x"7E",x"0E",x"80", -- 0x3220
		x"DD",x"77",x"0E",x"CB",x"78",x"C8",x"3F",x"C9", -- 0x3228
		x"DD",x"34",x"03",x"DD",x"5E",x"22",x"DD",x"56", -- 0x3230
		x"23",x"D5",x"FD",x"E1",x"FD",x"7E",x"0D",x"E6", -- 0x3238
		x"10",x"4F",x"DD",x"7E",x"0D",x"E6",x"EF",x"B1", -- 0x3240
		x"DD",x"77",x"0D",x"FD",x"7E",x"0F",x"DD",x"77", -- 0x3248
		x"0F",x"C3",x"E8",x"2A",x"CD",x"25",x"34",x"DD", -- 0x3250
		x"7E",x"08",x"E6",x"E0",x"20",x"19",x"DD",x"CB", -- 0x3258
		x"01",x"6E",x"C2",x"F7",x"43",x"DD",x"7E",x"12", -- 0x3260
		x"CD",x"F7",x"66",x"93",x"39",x"E4",x"3B",x"E4", -- 0x3268
		x"3B",x"39",x"3F",x"39",x"3F",x"A3",x"41",x"DD", -- 0x3270
		x"CB",x"02",x"66",x"CA",x"97",x"31",x"CD",x"F3", -- 0x3278
		x"31",x"F5",x"DD",x"35",x"16",x"CC",x"A2",x"32", -- 0x3280
		x"F1",x"D2",x"B4",x"31",x"DD",x"6E",x"1E",x"DD", -- 0x3288
		x"66",x"1F",x"23",x"35",x"CA",x"25",x"65",x"C3", -- 0x3290
		x"CB",x"66",x"CD",x"E8",x"2A",x"DD",x"36",x"00", -- 0x3298
		x"00",x"C9",x"DD",x"6E",x"10",x"DD",x"66",x"11", -- 0x32A0
		x"23",x"23",x"7E",x"B7",x"28",x"32",x"FE",x"FF", -- 0x32A8
		x"C2",x"CB",x"32",x"23",x"7E",x"E5",x"07",x"4F", -- 0x32B0
		x"06",x"00",x"21",x"8E",x"B1",x"09",x"7E",x"23", -- 0x32B8
		x"66",x"6F",x"DD",x"7E",x"08",x"E6",x"0F",x"4F", -- 0x32C0
		x"09",x"7E",x"E1",x"DD",x"77",x"16",x"23",x"CD", -- 0x32C8
		x"E5",x"32",x"23",x"DD",x"75",x"10",x"DD",x"74", -- 0x32D0
		x"11",x"CD",x"0A",x"42",x"DD",x"77",x"0C",x"C9", -- 0x32D8
		x"DD",x"36",x"16",x"7F",x"C9",x"7E",x"DD",x"CB", -- 0x32E0
		x"02",x"6E",x"28",x"35",x"FE",x"10",x"30",x"06", -- 0x32E8
		x"ED",x"44",x"E6",x"0F",x"18",x"2B",x"CB",x"5F", -- 0x32F0
		x"28",x"08",x"D6",x"10",x"EE",x"10",x"C6",x"10", -- 0x32F8
		x"18",x"1F",x"FE",x"28",x"30",x"1B",x"FE",x"20", -- 0x3300
		x"38",x"17",x"DD",x"CB",x"08",x"76",x"28",x"11", -- 0x3308
		x"4F",x"DD",x"7E",x"02",x"E6",x"0F",x"FE",x"03", -- 0x3310
		x"79",x"20",x"06",x"ED",x"44",x"E6",x"07",x"F6", -- 0x3318
		x"20",x"DD",x"77",x"19",x"C9",x"3A",x"99",x"E0", -- 0x3320
		x"B7",x"C0",x"DD",x"E5",x"FD",x"E1",x"CD",x"BE", -- 0x3328
		x"36",x"D0",x"CD",x"96",x"33",x"D8",x"B7",x"CC", -- 0x3330
		x"41",x"33",x"DD",x"CB",x"00",x"CE",x"C3",x"18", -- 0x3338
		x"36",x"3E",x"01",x"32",x"A5",x"E0",x"AF",x"01", -- 0x3340
		x"30",x"67",x"FF",x"C9",x"3A",x"99",x"E0",x"B7", -- 0x3348
		x"C0",x"3A",x"02",x"EC",x"FE",x"00",x"C0",x"21", -- 0x3350
		x"5C",x"37",x"DD",x"E5",x"FD",x"E1",x"CD",x"D4", -- 0x3358
		x"36",x"30",x"05",x"CD",x"96",x"33",x"30",x"0F", -- 0x3360
		x"21",x"60",x"37",x"DD",x"E5",x"FD",x"E1",x"CD", -- 0x3368
		x"11",x"37",x"D0",x"CD",x"96",x"33",x"D8",x"B7", -- 0x3370
		x"CC",x"41",x"33",x"C3",x"0D",x"36",x"3A",x"99", -- 0x3378
		x"E0",x"B7",x"C0",x"DD",x"E5",x"FD",x"E1",x"CD", -- 0x3380
		x"93",x"36",x"D0",x"CD",x"96",x"33",x"D8",x"B7", -- 0x3388
		x"CC",x"41",x"33",x"C3",x"1C",x"36",x"3A",x"A5", -- 0x3390
		x"E0",x"B7",x"20",x"1E",x"DD",x"7E",x"00",x"E6", -- 0x3398
		x"06",x"20",x"17",x"CD",x"19",x"34",x"C6",x"06", -- 0x33A0
		x"B8",x"38",x"0F",x"79",x"BC",x"38",x"0B",x"7B", -- 0x33A8
		x"BD",x"38",x"07",x"7D",x"C6",x"06",x"BA",x"3E", -- 0x33B0
		x"00",x"D0",x"3A",x"B4",x"E7",x"B7",x"20",x"40", -- 0x33B8
		x"3A",x"20",x"E1",x"6F",x"2F",x"E6",x"82",x"20", -- 0x33C0
		x"14",x"7D",x"E6",x"0C",x"20",x"0F",x"2A",x"2E", -- 0x33C8
		x"E1",x"CD",x"02",x"34",x"38",x"07",x"21",x"20", -- 0x33D0
		x"E1",x"CB",x"D6",x"18",x"1B",x"3A",x"30",x"E1", -- 0x33D8
		x"6F",x"2F",x"E6",x"82",x"20",x"1A",x"7D",x"E6", -- 0x33E0
		x"0C",x"20",x"15",x"2A",x"3E",x"E1",x"CD",x"02", -- 0x33E8
		x"34",x"38",x"0D",x"21",x"30",x"E1",x"CB",x"D6", -- 0x33F0
		x"DD",x"CB",x"00",x"CE",x"3E",x"01",x"B7",x"C9", -- 0x33F8
		x"37",x"C9",x"7D",x"C6",x"04",x"6F",x"7C",x"C6", -- 0x3400
		x"04",x"67",x"C6",x"05",x"B8",x"D8",x"79",x"BC", -- 0x3408
		x"D8",x"7B",x"BD",x"D8",x"7D",x"C6",x"04",x"BA", -- 0x3410
		x"C9",x"2A",x"0E",x"E1",x"7D",x"C6",x"0C",x"6F", -- 0x3418
		x"7C",x"C6",x"05",x"67",x"C9",x"06",x"03",x"FD", -- 0x3420
		x"21",x"60",x"E2",x"C5",x"FD",x"7E",x"00",x"CB", -- 0x3428
		x"47",x"28",x"0B",x"E6",x"0C",x"20",x"07",x"FD", -- 0x3430
		x"CB",x"01",x"46",x"CA",x"47",x"34",x"11",x"10", -- 0x3438
		x"00",x"FD",x"19",x"C1",x"10",x"E5",x"C9",x"DD", -- 0x3440
		x"7E",x"00",x"E6",x"C0",x"CA",x"DE",x"34",x"FE", -- 0x3448
		x"C0",x"CA",x"E8",x"34",x"FE",x"40",x"C2",x"3E", -- 0x3450
		x"34",x"DD",x"CB",x"01",x"76",x"C2",x"9B",x"35", -- 0x3458
		x"3A",x"02",x"EC",x"FE",x"00",x"C2",x"3E",x"34", -- 0x3460
		x"16",x"00",x"21",x"5C",x"37",x"CD",x"D4",x"36", -- 0x3468
		x"30",x"05",x"CD",x"27",x"36",x"30",x"0F",x"16", -- 0x3470
		x"01",x"21",x"60",x"37",x"CD",x"11",x"37",x"30", -- 0x3478
		x"BD",x"CD",x"27",x"36",x"38",x"B8",x"DD",x"34", -- 0x3480
		x"0A",x"21",x"64",x"37",x"CD",x"4E",x"37",x"DD", -- 0x3488
		x"4E",x"1D",x"09",x"DD",x"7E",x"0A",x"BE",x"D2", -- 0x3490
		x"AA",x"34",x"7E",x"DD",x"96",x"0A",x"FE",x"03", -- 0x3498
		x"D2",x"85",x"35",x"DD",x"CB",x"18",x"CE",x"C3", -- 0x34A0
		x"85",x"35",x"CD",x"76",x"36",x"FD",x"CB",x"01", -- 0x34A8
		x"C6",x"DD",x"CB",x"18",x"8E",x"21",x"00",x"00", -- 0x34B0
		x"22",x"70",x"E0",x"22",x"72",x"E0",x"22",x"76", -- 0x34B8
		x"E0",x"3A",x"07",x"EC",x"07",x"07",x"C6",x"02", -- 0x34C0
		x"4F",x"06",x"00",x"21",x"8C",x"7E",x"09",x"7E", -- 0x34C8
		x"32",x"74",x"E0",x"23",x"7E",x"32",x"75",x"E0", -- 0x34D0
		x"21",x"77",x"E0",x"C3",x"8E",x"35",x"DD",x"7E", -- 0x34D8
		x"01",x"E6",x"C0",x"FE",x"C0",x"CA",x"2B",x"35", -- 0x34E0
		x"CD",x"BE",x"36",x"D2",x"3E",x"34",x"CD",x"27", -- 0x34E8
		x"36",x"DA",x"3E",x"34",x"CD",x"76",x"36",x"FD", -- 0x34F0
		x"CB",x"01",x"C6",x"DD",x"7E",x"08",x"E6",x"E0", -- 0x34F8
		x"20",x"08",x"21",x"70",x"E1",x"7E",x"B7",x"28", -- 0x3500
		x"01",x"35",x"DD",x"7E",x"01",x"E6",x"C0",x"07", -- 0x3508
		x"07",x"07",x"4F",x"06",x"00",x"21",x"42",x"38", -- 0x3510
		x"09",x"7E",x"23",x"66",x"6F",x"DD",x"7E",x"1D", -- 0x3518
		x"E6",x"03",x"07",x"07",x"07",x"C6",x"07",x"4F", -- 0x3520
		x"09",x"18",x"63",x"CD",x"93",x"36",x"D2",x"3E", -- 0x3528
		x"34",x"CD",x"27",x"36",x"DA",x"3E",x"34",x"DD", -- 0x3530
		x"34",x"0A",x"DD",x"7E",x"08",x"E6",x"18",x"0F", -- 0x3538
		x"0F",x"4F",x"06",x"00",x"21",x"14",x"38",x"09", -- 0x3540
		x"7E",x"23",x"66",x"6F",x"CD",x"4E",x"37",x"DD", -- 0x3548
		x"4E",x"1D",x"09",x"DD",x"7E",x"0A",x"BE",x"30", -- 0x3550
		x"10",x"7E",x"DD",x"96",x"0A",x"FE",x"03",x"D2", -- 0x3558
		x"85",x"35",x"DD",x"CB",x"18",x"CE",x"C3",x"85", -- 0x3560
		x"35",x"FD",x"CB",x"01",x"C6",x"CD",x"76",x"36", -- 0x3568
		x"DD",x"CB",x"18",x"8E",x"DD",x"7E",x"1D",x"07", -- 0x3570
		x"07",x"07",x"C6",x"07",x"4F",x"06",x"00",x"21", -- 0x3578
		x"32",x"38",x"09",x"18",x"09",x"FD",x"CB",x"00", -- 0x3580
		x"D6",x"21",x"63",x"38",x"18",x"04",x"DD",x"CB", -- 0x3588
		x"00",x"CE",x"CD",x"D1",x"12",x"CD",x"55",x"2D", -- 0x3590
		x"C1",x"37",x"C9",x"21",x"D4",x"37",x"CD",x"6C", -- 0x3598
		x"37",x"30",x"05",x"CD",x"27",x"36",x"30",x"0F", -- 0x35A0
		x"21",x"D8",x"37",x"CD",x"A0",x"37",x"D2",x"3E", -- 0x35A8
		x"34",x"CD",x"27",x"36",x"DA",x"3E",x"34",x"DD", -- 0x35B0
		x"34",x"0A",x"21",x"DC",x"37",x"CD",x"4E",x"37", -- 0x35B8
		x"7E",x"23",x"66",x"6F",x"3A",x"03",x"E1",x"E6", -- 0x35C0
		x"18",x"0F",x"0F",x"0F",x"4F",x"09",x"DD",x"7E", -- 0x35C8
		x"0A",x"BE",x"D2",x"E6",x"35",x"7E",x"DD",x"96", -- 0x35D0
		x"0A",x"FE",x"03",x"D2",x"85",x"35",x"3E",x"01", -- 0x35D8
		x"32",x"F8",x"E9",x"C3",x"85",x"35",x"CD",x"76", -- 0x35E0
		x"36",x"FD",x"CB",x"01",x"C6",x"21",x"00",x"00", -- 0x35E8
		x"22",x"70",x"E0",x"22",x"72",x"E0",x"22",x"74", -- 0x35F0
		x"E0",x"22",x"76",x"E0",x"3A",x"03",x"E1",x"E6", -- 0x35F8
		x"18",x"C6",x"07",x"4F",x"06",x"00",x"21",x"F4", -- 0x3600
		x"37",x"09",x"C3",x"8E",x"35",x"C5",x"DD",x"CB", -- 0x3608
		x"18",x"8E",x"21",x"4F",x"38",x"C3",x"8E",x"35", -- 0x3610
		x"C5",x"C3",x"0A",x"35",x"C5",x"DD",x"CB",x"18", -- 0x3618
		x"8E",x"21",x"F1",x"52",x"C3",x"8E",x"35",x"79", -- 0x3620
		x"FD",x"BE",x"0F",x"D8",x"FD",x"7E",x"0F",x"C6", -- 0x3628
		x"05",x"B8",x"D8",x"FD",x"CB",x"00",x"6E",x"3A", -- 0x3630
		x"64",x"E1",x"28",x"09",x"07",x"3E",x"F3",x"38", -- 0x3638
		x"0B",x"D6",x"08",x"18",x"07",x"07",x"3E",x"02", -- 0x3640
		x"30",x"02",x"3E",x"07",x"FD",x"86",x"0E",x"4F", -- 0x3648
		x"7B",x"B9",x"D8",x"3A",x"64",x"E1",x"07",x"3E", -- 0x3650
		x"1C",x"38",x"0C",x"FD",x"CB",x"00",x"66",x"3E", -- 0x3658
		x"0C",x"28",x"0E",x"3E",x"22",x"18",x"0A",x"FD", -- 0x3660
		x"CB",x"00",x"66",x"3E",x"17",x"28",x"02",x"3E", -- 0x3668
		x"2A",x"FD",x"86",x"0E",x"BA",x"C9",x"21",x"4D", -- 0x3670
		x"E1",x"CD",x"8B",x"36",x"21",x"55",x"E1",x"C3", -- 0x3678
		x"8B",x"36",x"21",x"5D",x"E1",x"CD",x"8B",x"36", -- 0x3680
		x"21",x"65",x"E1",x"34",x"C0",x"23",x"34",x"C0", -- 0x3688
		x"23",x"34",x"C9",x"DD",x"7E",x"0D",x"E6",x"10", -- 0x3690
		x"DD",x"7E",x"0F",x"20",x"16",x"C6",x"03",x"D8", -- 0x3698
		x"47",x"C6",x"16",x"30",x"02",x"3E",x"FF",x"4F", -- 0x36A0
		x"DD",x"7E",x"0E",x"C6",x"08",x"57",x"C6",x"0F", -- 0x36A8
		x"5F",x"37",x"C9",x"C6",x"03",x"38",x"E9",x"C6", -- 0x36B0
		x"16",x"D0",x"06",x"00",x"18",x"E9",x"DD",x"7E", -- 0x36B8
		x"0D",x"E6",x"10",x"C0",x"DD",x"7E",x"0F",x"47", -- 0x36C0
		x"C6",x"0F",x"4F",x"DD",x"7E",x"0E",x"57",x"C6", -- 0x36C8
		x"0F",x"5F",x"37",x"C9",x"DD",x"5E",x"0D",x"DD", -- 0x36D0
		x"7E",x"0F",x"CB",x"63",x"28",x"13",x"FE",x"C0", -- 0x36D8
		x"DA",x"4C",x"37",x"06",x"00",x"7E",x"23",x"86", -- 0x36E0
		x"DD",x"86",x"0F",x"D2",x"4C",x"37",x"4F",x"18", -- 0x36E8
		x"0C",x"86",x"47",x"DA",x"4C",x"37",x"23",x"86", -- 0x36F0
		x"4F",x"30",x"02",x"0E",x"FF",x"23",x"DD",x"7E", -- 0x36F8
		x"0E",x"86",x"57",x"FE",x"F0",x"30",x"45",x"23", -- 0x3700
		x"86",x"5F",x"FE",x"F0",x"D8",x"1E",x"F0",x"37", -- 0x3708
		x"C9",x"3A",x"18",x"EC",x"5F",x"3A",x"1A",x"EC", -- 0x3710
		x"4F",x"79",x"CB",x"63",x"28",x"0F",x"FE",x"F1", -- 0x3718
		x"38",x"2A",x"06",x"00",x"7E",x"23",x"86",x"81", -- 0x3720
		x"30",x"22",x"4F",x"18",x"0B",x"86",x"38",x"1C", -- 0x3728
		x"47",x"23",x"86",x"4F",x"30",x"02",x"0E",x"FF", -- 0x3730
		x"23",x"3A",x"19",x"EC",x"86",x"FE",x"F0",x"30", -- 0x3738
		x"0B",x"57",x"23",x"86",x"FE",x"F0",x"5F",x"D8", -- 0x3740
		x"1E",x"EF",x"37",x"C9",x"B7",x"C9",x"3A",x"04", -- 0x3748
		x"C0",x"E6",x"60",x"0F",x"0F",x"0F",x"0F",x"4F", -- 0x3750
		x"06",x"00",x"09",x"C9",x"09",x"2C",x"0C",x"07", -- 0x3758
		x"02",x"06",x"08",x"30",x"19",x"1E",x"14",x"19", -- 0x3760
		x"0A",x"0F",x"0F",x"14",x"DD",x"5E",x"0D",x"DD", -- 0x3768
		x"7E",x"0F",x"CB",x"63",x"28",x"13",x"FE",x"80", -- 0x3770
		x"DA",x"D2",x"37",x"06",x"00",x"7E",x"23",x"86", -- 0x3778
		x"DD",x"86",x"0F",x"D2",x"D2",x"37",x"4F",x"18", -- 0x3780
		x"0C",x"86",x"47",x"DA",x"D2",x"37",x"23",x"86", -- 0x3788
		x"4F",x"30",x"02",x"0E",x"FF",x"23",x"DD",x"7E", -- 0x3790
		x"0E",x"86",x"57",x"23",x"86",x"5F",x"37",x"C9", -- 0x3798
		x"3A",x"51",x"EB",x"5F",x"3A",x"53",x"EB",x"4F", -- 0x37A0
		x"79",x"CB",x"63",x"28",x"0F",x"FE",x"F1",x"38", -- 0x37A8
		x"21",x"06",x"00",x"7E",x"23",x"86",x"81",x"30", -- 0x37B0
		x"19",x"4F",x"18",x"0B",x"86",x"38",x"13",x"47", -- 0x37B8
		x"23",x"86",x"4F",x"30",x"02",x"0E",x"FF",x"23", -- 0x37C0
		x"3A",x"52",x"EB",x"86",x"57",x"23",x"86",x"5F", -- 0x37C8
		x"37",x"C9",x"B7",x"C9",x"13",x"55",x"04",x"13", -- 0x37D0
		x"00",x"0F",x"0C",x"A6",x"F0",x"37",x"EC",x"37", -- 0x37D8
		x"E8",x"37",x"E4",x"37",x"28",x"2D",x"32",x"37", -- 0x37E0
		x"1E",x"23",x"28",x"2D",x"32",x"37",x"3C",x"42", -- 0x37E8
		x"46",x"4B",x"50",x"5A",x"00",x"00",x"00",x"02", -- 0x37F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03", -- 0x37F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04", -- 0x3800
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05", -- 0x3808
		x"00",x"00",x"00",x"00",x"1A",x"38",x"22",x"38", -- 0x3810
		x"2A",x"38",x"0A",x"0D",x"07",x"09",x"02",x"04", -- 0x3818
		x"04",x"06",x"0B",x"0D",x"08",x"0A",x"03",x"05", -- 0x3820
		x"05",x"07",x"0E",x"10",x"09",x"0B",x"04",x"06", -- 0x3828
		x"06",x"08",x"00",x"00",x"00",x"00",x"01",x"00", -- 0x3830
		x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"05", -- 0x3838
		x"00",x"00",x"4C",x"38",x"64",x"38",x"7C",x"38", -- 0x3840
		x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00", -- 0x3848
		x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"00", -- 0x3850
		x"00",x"00",x"05",x"00",x"00",x"00",x"00",x"00", -- 0x3858
		x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3860
		x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00", -- 0x3868
		x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3870
		x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3878
		x"00",x"01",x"05",x"00",x"00",x"00",x"00",x"00", -- 0x3880
		x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3888
		x"00",x"02",x"00",x"00",x"DD",x"5E",x"0F",x"1C", -- 0x3890
		x"2A",x"0E",x"E1",x"7C",x"C6",x"0C",x"BB",x"D8", -- 0x3898
		x"D6",x"08",x"BB",x"3F",x"D8",x"7D",x"C6",x"08", -- 0x38A0
		x"6F",x"DD",x"7E",x"0E",x"C6",x"08",x"BD",x"D8", -- 0x38A8
		x"4F",x"7D",x"C6",x"10",x"B9",x"C9",x"FD",x"21", -- 0x38B0
		x"20",x"E1",x"CD",x"C2",x"38",x"D0",x"FD",x"21", -- 0x38B8
		x"30",x"E1",x"FD",x"7E",x"00",x"5F",x"2F",x"E6", -- 0x38C0
		x"82",x"37",x"C0",x"7B",x"E6",x"3C",x"37",x"C0", -- 0x38C8
		x"DD",x"5E",x"0F",x"1C",x"FD",x"6E",x"0E",x"FD", -- 0x38D0
		x"66",x"0F",x"7C",x"C6",x"0C",x"BB",x"D8",x"D6", -- 0x38D8
		x"08",x"BB",x"3F",x"D8",x"7D",x"C6",x"04",x"6F", -- 0x38E0
		x"DD",x"7E",x"0E",x"C6",x"08",x"BD",x"D8",x"4F", -- 0x38E8
		x"7D",x"C6",x"08",x"B9",x"D8",x"FD",x"CB",x"00", -- 0x38F0
		x"D6",x"C9",x"CD",x"D4",x"56",x"E6",x"3F",x"4F", -- 0x38F8
		x"CB",x"76",x"06",x"08",x"28",x"02",x"06",x"A8", -- 0x3900
		x"80",x"DD",x"77",x"0E",x"DD",x"36",x"0C",x"20", -- 0x3908
		x"DD",x"36",x"19",x"0C",x"DD",x"36",x"0F",x"FF", -- 0x3910
		x"DD",x"36",x"14",x"06",x"DD",x"36",x"02",x"02", -- 0x3918
		x"DD",x"34",x"03",x"C9",x"01",x"C0",x"8B",x"CD", -- 0x3920
		x"85",x"3B",x"AF",x"DD",x"77",x"17",x"DD",x"77", -- 0x3928
		x"14",x"DD",x"36",x"09",x"02",x"2A",x"0E",x"E1", -- 0x3930
		x"01",x"08",x"00",x"09",x"DD",x"7E",x"0F",x"94", -- 0x3938
		x"DC",x"90",x"39",x"0F",x"0F",x"0F",x"0F",x"E6", -- 0x3940
		x"0F",x"67",x"0E",x"00",x"DD",x"7E",x"0E",x"95", -- 0x3948
		x"D4",x"8E",x"39",x"0F",x"0F",x"0F",x"E6",x"1F", -- 0x3950
		x"6F",x"BC",x"20",x"04",x"0E",x"04",x"18",x"03", -- 0x3958
		x"30",x"01",x"0C",x"DD",x"7E",x"01",x"E6",x"C0", -- 0x3960
		x"B1",x"DD",x"77",x"01",x"DD",x"7E",x"19",x"FE", -- 0x3968
		x"30",x"38",x"04",x"E6",x"7C",x"18",x"0D",x"E6", -- 0x3970
		x"3C",x"FE",x"10",x"30",x"05",x"07",x"C6",x"30", -- 0x3978
		x"18",x"02",x"C6",x"20",x"DD",x"77",x"19",x"CD", -- 0x3980
		x"10",x"42",x"DD",x"34",x"03",x"C9",x"0E",x"02", -- 0x3988
		x"ED",x"44",x"C9",x"CD",x"EC",x"50",x"DD",x"56", -- 0x3990
		x"02",x"CB",x"52",x"20",x"5C",x"CD",x"CB",x"3A", -- 0x3998
		x"D8",x"DD",x"CB",x"02",x"6E",x"C2",x"1C",x"3A", -- 0x39A0
		x"DD",x"CB",x"0D",x"66",x"C2",x"E8",x"2A",x"DD", -- 0x39A8
		x"5E",x"02",x"16",x"14",x"CB",x"43",x"28",x"02", -- 0x39B0
		x"16",x"F8",x"3A",x"0F",x"E1",x"E6",x"F8",x"82", -- 0x39B8
		x"4F",x"DD",x"7E",x"0F",x"E6",x"F8",x"B9",x"28", -- 0x39C0
		x"26",x"CB",x"43",x"28",x"01",x"3F",x"DA",x"EF", -- 0x39C8
		x"39",x"3A",x"0E",x"E1",x"C6",x"08",x"DD",x"96", -- 0x39D0
		x"0E",x"DC",x"90",x"39",x"FE",x"30",x"D2",x"E8", -- 0x39D8
		x"2A",x"3A",x"0F",x"E1",x"DD",x"96",x"0F",x"DC", -- 0x39E0
		x"90",x"39",x"FE",x"58",x"D2",x"E8",x"2A",x"DD", -- 0x39E8
		x"CB",x"02",x"D6",x"CD",x"2F",x"3A",x"C3",x"E8", -- 0x39F0
		x"2A",x"CD",x"AA",x"3A",x"D8",x"DD",x"35",x"16", -- 0x39F8
		x"C2",x"E8",x"2A",x"CD",x"73",x"3A",x"D2",x"E8", -- 0x3A00
		x"2A",x"DD",x"7E",x"02",x"E6",x"FB",x"EE",x"09", -- 0x3A08
		x"F6",x"20",x"DD",x"77",x"02",x"DD",x"36",x"16", -- 0x3A10
		x"20",x"C3",x"E8",x"2A",x"DD",x"35",x"16",x"C2", -- 0x3A18
		x"E8",x"2A",x"CD",x"38",x"4E",x"DA",x"E8",x"2A", -- 0x3A20
		x"DD",x"36",x"16",x"FF",x"C3",x"E8",x"2A",x"16", -- 0x3A28
		x"00",x"21",x"9F",x"79",x"DD",x"7E",x"01",x"CB", -- 0x3A30
		x"57",x"20",x"0D",x"CB",x"4F",x"28",x"02",x"16", -- 0x3A38
		x"10",x"E6",x"01",x"3C",x"07",x"4F",x"18",x"0E", -- 0x3A40
		x"3A",x"0E",x"E1",x"C6",x"08",x"DD",x"BE",x"0E", -- 0x3A48
		x"30",x"02",x"16",x"10",x"0E",x"00",x"06",x"00", -- 0x3A50
		x"09",x"7E",x"23",x"66",x"6F",x"7E",x"DD",x"77", -- 0x3A58
		x"16",x"23",x"23",x"DD",x"75",x"1E",x"DD",x"74", -- 0x3A60
		x"1F",x"DD",x"7E",x"01",x"E6",x"EF",x"B2",x"DD", -- 0x3A68
		x"77",x"01",x"C9",x"DD",x"6E",x"1E",x"DD",x"66", -- 0x3A70
		x"1F",x"23",x"23",x"7E",x"B7",x"28",x"29",x"DD", -- 0x3A78
		x"77",x"16",x"23",x"56",x"23",x"DD",x"75",x"1E", -- 0x3A80
		x"DD",x"74",x"1F",x"DD",x"CB",x"02",x"5E",x"28", -- 0x3A88
		x"0C",x"7A",x"C6",x"04",x"57",x"E6",x"07",x"20", -- 0x3A90
		x"04",x"7A",x"D6",x"08",x"57",x"DD",x"72",x"19", -- 0x3A98
		x"CD",x"10",x"42",x"DD",x"77",x"0C",x"B7",x"C9", -- 0x3AA0
		x"37",x"C9",x"DD",x"6E",x"1E",x"DD",x"66",x"1F", -- 0x3AA8
		x"4E",x"23",x"46",x"DD",x"CB",x"02",x"5E",x"28", -- 0x3AB0
		x"04",x"79",x"ED",x"44",x"4F",x"DD",x"CB",x"01", -- 0x3AB8
		x"66",x"CA",x"FB",x"3A",x"78",x"ED",x"44",x"47", -- 0x3AC0
		x"C3",x"FB",x"3A",x"06",x"00",x"0E",x"FE",x"DD", -- 0x3AC8
		x"56",x"01",x"CB",x"52",x"20",x"1A",x"04",x"CB", -- 0x3AD0
		x"42",x"20",x"0D",x"DD",x"7E",x"17",x"EE",x"20", -- 0x3AD8
		x"DD",x"77",x"17",x"E6",x"20",x"20",x"01",x"05", -- 0x3AE0
		x"CB",x"4A",x"28",x"04",x"78",x"ED",x"44",x"47", -- 0x3AE8
		x"DD",x"CB",x"02",x"46",x"CA",x"FB",x"3A",x"79", -- 0x3AF0
		x"ED",x"44",x"4F",x"78",x"B7",x"CA",x"16",x"3B", -- 0x3AF8
		x"CB",x"7F",x"20",x"0A",x"DD",x"86",x"0E",x"DD", -- 0x3B00
		x"77",x"0E",x"38",x"3C",x"18",x"08",x"DD",x"86", -- 0x3B08
		x"0E",x"DD",x"77",x"0E",x"30",x"32",x"79",x"B7", -- 0x3B10
		x"C8",x"CB",x"7F",x"20",x"12",x"DD",x"86",x"0F", -- 0x3B18
		x"DD",x"77",x"0F",x"D0",x"DD",x"CB",x"0D",x"66", -- 0x3B20
		x"28",x"1E",x"DD",x"CB",x"0D",x"A6",x"C9",x"DD", -- 0x3B28
		x"86",x"0F",x"DD",x"77",x"0F",x"3F",x"DD",x"CB", -- 0x3B30
		x"0D",x"66",x"38",x"03",x"C8",x"18",x"06",x"20", -- 0x3B38
		x"07",x"DD",x"CB",x"0D",x"E6",x"FE",x"F1",x"D0", -- 0x3B40
		x"CD",x"6A",x"3B",x"18",x"04",x"CD",x"56",x"3B", -- 0x3B48
		x"D0",x"CD",x"CB",x"66",x"37",x"C9",x"DD",x"CB", -- 0x3B50
		x"0D",x"66",x"28",x"07",x"DD",x"7E",x"0F",x"FE", -- 0x3B58
		x"F1",x"38",x"07",x"DD",x"7E",x"0E",x"FE",x"F2", -- 0x3B60
		x"3F",x"D0",x"DD",x"7E",x"08",x"E6",x"E0",x"20", -- 0x3B68
		x"0F",x"DD",x"7E",x"00",x"E6",x"C0",x"20",x"08", -- 0x3B70
		x"21",x"70",x"E1",x"7E",x"B7",x"28",x"01",x"35", -- 0x3B78
		x"37",x"C9",x"01",x"C0",x"83",x"DD",x"7E",x"02", -- 0x3B80
		x"A0",x"DD",x"77",x"02",x"DD",x"7E",x"01",x"A1", -- 0x3B88
		x"DD",x"77",x"01",x"C9",x"CD",x"D4",x"56",x"E6", -- 0x3B90
		x"7F",x"C6",x"30",x"DD",x"77",x"0E",x"DD",x"36", -- 0x3B98
		x"19",x"20",x"DD",x"36",x"0C",x"20",x"C3",x"14", -- 0x3BA0
		x"39",x"DD",x"CB",x"02",x"DE",x"01",x"C0",x"8B", -- 0x3BA8
		x"18",x"03",x"01",x"C0",x"83",x"CD",x"85",x"3B", -- 0x3BB0
		x"AF",x"DD",x"77",x"13",x"DD",x"77",x"14",x"DD", -- 0x3BB8
		x"77",x"15",x"3E",x"02",x"DD",x"77",x"09",x"DD", -- 0x3BC0
		x"7E",x"19",x"FE",x"10",x"38",x"0A",x"FE",x"30", -- 0x3BC8
		x"38",x"0E",x"D6",x"30",x"E6",x"18",x"18",x"03", -- 0x3BD0
		x"E6",x"0C",x"07",x"C6",x"10",x"DD",x"77",x"19", -- 0x3BD8
		x"DD",x"34",x"03",x"C9",x"CD",x"EC",x"50",x"DD", -- 0x3BE0
		x"CB",x"02",x"56",x"20",x"73",x"DD",x"CB",x"02", -- 0x3BE8
		x"76",x"20",x"5F",x"3A",x"0F",x"E1",x"4F",x"CD", -- 0x3BF0
		x"09",x"62",x"AF",x"47",x"ED",x"42",x"7C",x"B7", -- 0x3BF8
		x"20",x"50",x"7D",x"FE",x"58",x"16",x"80",x"5F", -- 0x3C00
		x"30",x"48",x"3A",x"0E",x"E1",x"C6",x"08",x"DD", -- 0x3C08
		x"96",x"0E",x"30",x"02",x"ED",x"44",x"57",x"1E", -- 0x3C10
		x"80",x"FE",x"40",x"30",x"35",x"3A",x"0E",x"E1", -- 0x3C18
		x"C6",x"08",x"DD",x"BE",x"0E",x"01",x"04",x"27", -- 0x3C20
		x"16",x"27",x"30",x"05",x"01",x"0C",x"21",x"16", -- 0x3C28
		x"21",x"DD",x"7E",x"02",x"E6",x"03",x"B1",x"DD", -- 0x3C30
		x"77",x"02",x"DD",x"70",x"0C",x"DD",x"72",x"19", -- 0x3C38
		x"AF",x"DD",x"77",x"15",x"21",x"CC",x"7B",x"7E", -- 0x3C40
		x"DD",x"77",x"16",x"23",x"DD",x"75",x"1E",x"DD", -- 0x3C48
		x"74",x"1F",x"CD",x"FF",x"3C",x"D8",x"C3",x"E8", -- 0x3C50
		x"2A",x"CD",x"4D",x"3B",x"D8",x"C3",x"E8",x"2A", -- 0x3C58
		x"CD",x"C9",x"3C",x"D8",x"DD",x"35",x"16",x"C2", -- 0x3C60
		x"E8",x"2A",x"DD",x"34",x"15",x"DD",x"7E",x"15", -- 0x3C68
		x"FE",x"09",x"28",x"04",x"FE",x"0D",x"20",x"2E", -- 0x3C70
		x"DD",x"56",x"19",x"7A",x"E6",x"07",x"DD",x"CB", -- 0x3C78
		x"02",x"5E",x"28",x"0D",x"FE",x"07",x"38",x"06", -- 0x3C80
		x"7A",x"E6",x"30",x"57",x"18",x"0F",x"14",x"18", -- 0x3C88
		x"0C",x"B7",x"20",x"08",x"7A",x"E6",x"30",x"F6", -- 0x3C90
		x"07",x"57",x"18",x"01",x"15",x"DD",x"72",x"19", -- 0x3C98
		x"CD",x"10",x"42",x"DD",x"77",x"0C",x"CD",x"B3", -- 0x3CA0
		x"3C",x"C2",x"E8",x"2A",x"DD",x"36",x"16",x"FF", -- 0x3CA8
		x"C3",x"E8",x"2A",x"DD",x"6E",x"1E",x"DD",x"66", -- 0x3CB0
		x"1F",x"23",x"23",x"7E",x"B7",x"C8",x"DD",x"77", -- 0x3CB8
		x"16",x"23",x"DD",x"75",x"1E",x"DD",x"74",x"1F", -- 0x3CC0
		x"C9",x"DD",x"6E",x"1E",x"DD",x"66",x"1F",x"4E", -- 0x3CC8
		x"23",x"46",x"DD",x"CB",x"02",x"5E",x"CA",x"FB", -- 0x3CD0
		x"3A",x"78",x"ED",x"44",x"47",x"C3",x"FB",x"3A", -- 0x3CD8
		x"09",x"4E",x"23",x"46",x"C5",x"CB",x"79",x"06", -- 0x3CE0
		x"00",x"28",x"01",x"05",x"CD",x"F8",x"3C",x"C1", -- 0x3CE8
		x"DD",x"7E",x"0E",x"80",x"DD",x"77",x"0E",x"C9", -- 0x3CF0
		x"CD",x"09",x"62",x"09",x"C3",x"C8",x"50",x"21", -- 0x3CF8
		x"24",x"7C",x"DD",x"CB",x"02",x"76",x"28",x"03", -- 0x3D00
		x"21",x"2C",x"7C",x"DD",x"7E",x"02",x"E6",x"03", -- 0x3D08
		x"07",x"4F",x"06",x"00",x"09",x"4E",x"23",x"46", -- 0x3D10
		x"C3",x"FB",x"3A",x"CD",x"D4",x"56",x"E6",x"7F", -- 0x3D18
		x"C6",x"50",x"DD",x"77",x"0E",x"DD",x"36",x"19", -- 0x3D20
		x"20",x"DD",x"36",x"0C",x"20",x"C3",x"14",x"39", -- 0x3D28
		x"CD",x"D4",x"56",x"0F",x"0F",x"E6",x"03",x"CD", -- 0x3D30
		x"F7",x"66",x"42",x"3D",x"7E",x"3D",x"97",x"3D", -- 0x3D38
		x"BE",x"3D",x"CD",x"E5",x"3D",x"DD",x"36",x"0E", -- 0x3D40
		x"01",x"DD",x"36",x"19",x"08",x"CD",x"10",x"42", -- 0x3D48
		x"DD",x"77",x"0C",x"DD",x"36",x"14",x"00",x"0E", -- 0x3D50
		x"02",x"18",x"0E",x"CD",x"D4",x"56",x"E6",x"1F", -- 0x3D58
		x"C6",x"02",x"DD",x"77",x"17",x"DD",x"CB",x"01", -- 0x3D60
		x"DE",x"DD",x"7E",x"02",x"E6",x"80",x"B1",x"DD", -- 0x3D68
		x"77",x"02",x"DD",x"36",x"09",x"02",x"AF",x"DD", -- 0x3D70
		x"77",x"13",x"DD",x"34",x"03",x"C9",x"CD",x"FC", -- 0x3D78
		x"3D",x"DD",x"36",x"19",x"00",x"DD",x"36",x"0E", -- 0x3D80
		x"EF",x"CD",x"10",x"42",x"DD",x"77",x"0C",x"DD", -- 0x3D88
		x"36",x"14",x"03",x"0E",x"03",x"18",x"D2",x"CD", -- 0x3D90
		x"1A",x"3E",x"06",x"80",x"3A",x"03",x"E1",x"BE", -- 0x3D98
		x"38",x"02",x"06",x"58",x"CD",x"09",x"3E",x"DD", -- 0x3DA0
		x"36",x"19",x"04",x"DD",x"36",x"0E",x"EF",x"CD", -- 0x3DA8
		x"10",x"42",x"DD",x"77",x"0C",x"DD",x"36",x"14", -- 0x3DB0
		x"05",x"0E",x"01",x"C3",x"5B",x"3D",x"CD",x"1A", -- 0x3DB8
		x"3E",x"06",x"90",x"3A",x"03",x"E1",x"BE",x"38", -- 0x3DC0
		x"02",x"06",x"68",x"CD",x"09",x"3E",x"DD",x"36", -- 0x3DC8
		x"19",x"04",x"DD",x"36",x"0E",x"EF",x"CD",x"10", -- 0x3DD0
		x"42",x"DD",x"77",x"0C",x"DD",x"36",x"14",x"05", -- 0x3DD8
		x"0E",x"01",x"C3",x"69",x"3D",x"CD",x"1A",x"3E", -- 0x3DE0
		x"06",x"E0",x"3A",x"03",x"E1",x"BE",x"38",x"02", -- 0x3DE8
		x"06",x"90",x"3A",x"0C",x"E0",x"E6",x"1F",x"80", -- 0x3DF0
		x"DD",x"77",x"0F",x"C9",x"CD",x"1A",x"3E",x"06", -- 0x3DF8
		x"50",x"3A",x"03",x"E1",x"BE",x"30",x"02",x"06", -- 0x3E00
		x"80",x"3A",x"0C",x"E0",x"E6",x"1F",x"4F",x"3A", -- 0x3E08
		x"0E",x"E1",x"E6",x"1F",x"81",x"80",x"DD",x"77", -- 0x3E10
		x"0F",x"C9",x"21",x"C2",x"3E",x"3A",x"04",x"C0", -- 0x3E18
		x"E6",x"60",x"07",x"07",x"07",x"4F",x"06",x"00", -- 0x3E20
		x"09",x"C9",x"CD",x"D4",x"56",x"3A",x"0C",x"E0", -- 0x3E28
		x"86",x"0F",x"0F",x"E6",x"03",x"CD",x"F7",x"66", -- 0x3E30
		x"40",x"3E",x"67",x"3E",x"8E",x"3E",x"A8",x"3E", -- 0x3E38
		x"CD",x"1A",x"3E",x"06",x"90",x"3A",x"03",x"E1", -- 0x3E40
		x"BE",x"38",x"02",x"06",x"68",x"CD",x"09",x"3E", -- 0x3E48
		x"DD",x"36",x"0E",x"01",x"DD",x"36",x"19",x"0C", -- 0x3E50
		x"CD",x"10",x"42",x"DD",x"77",x"0C",x"DD",x"36", -- 0x3E58
		x"14",x"04",x"0E",x"08",x"C3",x"69",x"3D",x"CD", -- 0x3E60
		x"1A",x"3E",x"06",x"80",x"3A",x"03",x"E1",x"BE", -- 0x3E68
		x"38",x"02",x"06",x"58",x"CD",x"09",x"3E",x"DD", -- 0x3E70
		x"36",x"0E",x"01",x"DD",x"36",x"19",x"0C",x"CD", -- 0x3E78
		x"10",x"42",x"DD",x"77",x"0C",x"DD",x"36",x"14", -- 0x3E80
		x"04",x"0E",x"08",x"C3",x"5B",x"3D",x"CD",x"FC", -- 0x3E88
		x"3D",x"DD",x"36",x"0E",x"01",x"DD",x"36",x"19", -- 0x3E90
		x"00",x"CD",x"10",x"42",x"DD",x"77",x"0C",x"DD", -- 0x3E98
		x"36",x"14",x"02",x"0E",x"0B",x"C3",x"69",x"3D", -- 0x3EA0
		x"CD",x"E5",x"3D",x"DD",x"36",x"0E",x"EF",x"DD", -- 0x3EA8
		x"36",x"19",x"08",x"CD",x"10",x"42",x"DD",x"77", -- 0x3EB0
		x"0C",x"DD",x"36",x"14",x"01",x"0E",x"0A",x"C3", -- 0x3EB8
		x"69",x"3D",x"02",x"0D",x"20",x"20",x"CD",x"D4", -- 0x3EC0
		x"56",x"7E",x"E6",x"03",x"CA",x"42",x"3D",x"3D", -- 0x3EC8
		x"CA",x"BE",x"3D",x"3D",x"CA",x"7E",x"3D",x"DD", -- 0x3ED0
		x"7E",x"1A",x"FE",x"01",x"C2",x"97",x"3D",x"DD", -- 0x3ED8
		x"CB",x"01",x"E6",x"C3",x"97",x"3D",x"CD",x"D4", -- 0x3EE0
		x"56",x"7E",x"E6",x"03",x"CA",x"A8",x"3E",x"3D", -- 0x3EE8
		x"CA",x"40",x"3E",x"3D",x"CA",x"8E",x"3E",x"DD", -- 0x3EF0
		x"7E",x"1A",x"FE",x"01",x"C2",x"67",x"3E",x"DD", -- 0x3EF8
		x"CB",x"01",x"E6",x"C3",x"67",x"3E",x"DD",x"7E", -- 0x3F00
		x"02",x"E6",x"83",x"DD",x"77",x"02",x"DD",x"36", -- 0x3F08
		x"09",x"02",x"DD",x"7E",x"01",x"E6",x"C8",x"DD", -- 0x3F10
		x"77",x"01",x"DD",x"7E",x"19",x"FE",x"10",x"38", -- 0x3F18
		x"08",x"D6",x"10",x"E6",x"18",x"0F",x"DD",x"77", -- 0x3F20
		x"19",x"DD",x"34",x"03",x"C9",x"DD",x"7E",x"02", -- 0x3F28
		x"E6",x"83",x"F6",x"08",x"DD",x"77",x"02",x"18", -- 0x3F30
		x"D5",x"CD",x"EC",x"50",x"DD",x"CB",x"02",x"56", -- 0x3F38
		x"C2",x"87",x"40",x"DD",x"CB",x"01",x"56",x"C2", -- 0x3F40
		x"22",x"40",x"0E",x"00",x"DD",x"CB",x"0D",x"66", -- 0x3F48
		x"3A",x"0F",x"E1",x"20",x"0A",x"DD",x"96",x"0F", -- 0x3F50
		x"30",x"0C",x"0C",x"ED",x"44",x"18",x"07",x"5F", -- 0x3F58
		x"DD",x"7E",x"0F",x"ED",x"44",x"83",x"5F",x"3A", -- 0x3F60
		x"0E",x"E1",x"C6",x"08",x"DD",x"96",x"0E",x"30", -- 0x3F68
		x"04",x"ED",x"44",x"CB",x"C9",x"57",x"BB",x"30", -- 0x3F70
		x"01",x"7B",x"0F",x"0F",x"0F",x"E6",x"1F",x"5F", -- 0x3F78
		x"21",x"3E",x"7C",x"DD",x"CB",x"02",x"5E",x"28", -- 0x3F80
		x"03",x"21",x"42",x"7C",x"DD",x"7E",x"02",x"E6", -- 0x3F88
		x"03",x"06",x"00",x"09",x"BE",x"28",x"03",x"AF", -- 0x3F90
		x"18",x"18",x"7B",x"DD",x"CB",x"01",x"56",x"20", -- 0x3F98
		x"0B",x"FE",x"05",x"30",x"03",x"AF",x"18",x"0A", -- 0x3FA0
		x"FE",x"0F",x"38",x"02",x"3E",x"0F",x"D6",x"05", -- 0x3FA8
		x"E6",x"FE",x"21",x"9C",x"87",x"4F",x"06",x"00", -- 0x3FB0
		x"09",x"7E",x"23",x"66",x"6F",x"DD",x"7E",x"02", -- 0x3FB8
		x"E6",x"03",x"E2",x"C7",x"3F",x"EE",x"03",x"DD", -- 0x3FC0
		x"CB",x"02",x"5E",x"28",x"08",x"DD",x"CB",x"02", -- 0x3FC8
		x"4E",x"20",x"02",x"EE",x"02",x"FE",x"02",x"38", -- 0x3FD0
		x"02",x"D6",x"02",x"CD",x"09",x"41",x"7E",x"23", -- 0x3FD8
		x"66",x"6F",x"7E",x"DD",x"77",x"16",x"23",x"CD", -- 0x3FE0
		x"63",x"40",x"CD",x"10",x"42",x"DD",x"77",x"0C", -- 0x3FE8
		x"23",x"DD",x"75",x"1E",x"DD",x"74",x"1F",x"DD", -- 0x3FF0
		x"CB",x"02",x"D6",x"DD",x"56",x"19",x"DD",x"5E"  -- 0x3FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
