-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_M4 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_M4 is


	type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"01",x"7A",x"E6",x"03",x"28",x"04",x"CB",x"CB", -- 0x0000
		x"18",x"08",x"CB",x"8B",x"CB",x"43",x"20",x"0B", -- 0x0008
		x"CB",x"C3",x"7A",x"E6",x"0C",x"DD",x"77",x"1B", -- 0x0010
		x"DD",x"73",x"01",x"CD",x"3A",x"40",x"D2",x"E8", -- 0x0018
		x"2A",x"C9",x"DD",x"7E",x"19",x"FE",x"08",x"C2", -- 0x0020
		x"4A",x"3F",x"3A",x"C7",x"E0",x"B7",x"C2",x"4A", -- 0x0028
		x"3F",x"CD",x"38",x"4E",x"D2",x"4A",x"3F",x"C3", -- 0x0030
		x"E8",x"2A",x"4E",x"23",x"46",x"DD",x"56",x"02", -- 0x0038
		x"CB",x"5A",x"20",x"0B",x"CB",x"42",x"C2",x"FB", -- 0x0040
		x"3A",x"79",x"ED",x"44",x"4F",x"18",x"0D",x"7A", -- 0x0048
		x"E6",x"03",x"EA",x"5C",x"40",x"79",x"ED",x"44", -- 0x0050
		x"4F",x"C3",x"FB",x"3A",x"78",x"ED",x"44",x"47", -- 0x0058
		x"C3",x"FB",x"3A",x"7E",x"DD",x"CB",x"02",x"5E", -- 0x0060
		x"20",x"0A",x"DD",x"CB",x"02",x"46",x"20",x"13", -- 0x0068
		x"C6",x"08",x"18",x"0D",x"DD",x"7E",x"02",x"E6", -- 0x0070
		x"03",x"7E",x"EA",x"7F",x"40",x"C6",x"08",x"ED", -- 0x0078
		x"44",x"E6",x"0F",x"DD",x"77",x"19",x"C9",x"DD", -- 0x0080
		x"6E",x"1E",x"DD",x"66",x"1F",x"E5",x"CD",x"3A", -- 0x0088
		x"40",x"E1",x"D8",x"23",x"23",x"3A",x"C7",x"E0", -- 0x0090
		x"B7",x"C2",x"E8",x"2A",x"DD",x"35",x"16",x"C2", -- 0x0098
		x"E8",x"2A",x"7E",x"B7",x"CA",x"C6",x"40",x"DD", -- 0x00A0
		x"77",x"16",x"23",x"CD",x"63",x"40",x"E6",x"03", -- 0x00A8
		x"28",x"04",x"DD",x"CB",x"01",x"CE",x"CD",x"10", -- 0x00B0
		x"42",x"DD",x"77",x"0C",x"23",x"DD",x"75",x"1E", -- 0x00B8
		x"DD",x"74",x"1F",x"C3",x"E8",x"2A",x"DD",x"7E", -- 0x00C0
		x"19",x"5F",x"DD",x"BE",x"1B",x"20",x"08",x"DD", -- 0x00C8
		x"CB",x"01",x"86",x"DD",x"CB",x"01",x"D6",x"7B", -- 0x00D0
		x"E6",x"0C",x"E2",x"DF",x"40",x"EE",x"0C",x"0F", -- 0x00D8
		x"0F",x"5F",x"DD",x"7E",x"02",x"E6",x"F8",x"B3", -- 0x00E0
		x"DD",x"77",x"02",x"DD",x"CB",x"01",x"8E",x"C3", -- 0x00E8
		x"E8",x"2A",x"CD",x"0F",x"41",x"CD",x"E4",x"3C", -- 0x00F0
		x"DD",x"35",x"17",x"C2",x"59",x"3C",x"DD",x"CB", -- 0x00F8
		x"01",x"9E",x"C3",x"59",x"3C",x"DD",x"7E",x"15", -- 0x0100
		x"07",x"07",x"4F",x"06",x"00",x"09",x"C9",x"DD", -- 0x0108
		x"46",x"09",x"0E",x"00",x"DD",x"7E",x"02",x"E6", -- 0x0110
		x"03",x"C8",x"57",x"78",x"ED",x"44",x"47",x"15", -- 0x0118
		x"C8",x"48",x"06",x"00",x"15",x"C8",x"DD",x"4E", -- 0x0120
		x"09",x"C9",x"CD",x"D4",x"56",x"E6",x"1F",x"C6", -- 0x0128
		x"80",x"DD",x"77",x"0F",x"DD",x"36",x"02",x"00", -- 0x0130
		x"CB",x"5F",x"11",x"30",x"28",x"01",x"04",x"01", -- 0x0138
		x"28",x"06",x"01",x"05",x"EF",x"11",x"10",x"18", -- 0x0140
		x"DD",x"70",x"0E",x"DD",x"71",x"14",x"DD",x"73", -- 0x0148
		x"0C",x"DD",x"72",x"19",x"DD",x"6E",x"10",x"DD", -- 0x0150
		x"66",x"11",x"23",x"23",x"7E",x"FE",x"03",x"28", -- 0x0158
		x"04",x"DD",x"CB",x"02",x"DE",x"DD",x"7E",x"02", -- 0x0160
		x"B1",x"E6",x"FB",x"DD",x"77",x"02",x"DD",x"34", -- 0x0168
		x"03",x"C9",x"DD",x"CB",x"02",x"A6",x"DD",x"36", -- 0x0170
		x"14",x"04",x"DD",x"36",x"15",x"01",x"DD",x"7E", -- 0x0178
		x"19",x"FE",x"10",x"38",x"0E",x"FE",x"30",x"38", -- 0x0180
		x"12",x"E6",x"7C",x"D6",x"30",x"EE",x"10",x"C6", -- 0x0188
		x"10",x"18",x"05",x"E6",x"0C",x"07",x"C6",x"10", -- 0x0190
		x"DD",x"77",x"19",x"DD",x"36",x"09",x"02",x"DD", -- 0x0198
		x"34",x"03",x"C9",x"DD",x"35",x"15",x"20",x"34", -- 0x01A0
		x"DD",x"7E",x"14",x"DD",x"77",x"15",x"DD",x"46", -- 0x01A8
		x"19",x"78",x"E6",x"07",x"DD",x"CB",x"02",x"66", -- 0x01B0
		x"20",x"0D",x"FE",x"07",x"38",x"06",x"78",x"E6", -- 0x01B8
		x"38",x"47",x"18",x"0F",x"04",x"18",x"0C",x"B7", -- 0x01C0
		x"20",x"08",x"78",x"E6",x"38",x"F6",x"07",x"47", -- 0x01C8
		x"18",x"01",x"05",x"DD",x"70",x"19",x"CD",x"10", -- 0x01D0
		x"42",x"DD",x"77",x"0C",x"DD",x"46",x"09",x"58", -- 0x01D8
		x"0E",x"00",x"DD",x"7E",x"02",x"E6",x"03",x"57", -- 0x01E0
		x"28",x"0E",x"78",x"ED",x"44",x"47",x"15",x"28", -- 0x01E8
		x"07",x"48",x"06",x"00",x"15",x"28",x"01",x"4B", -- 0x01F0
		x"CD",x"FB",x"3A",x"D8",x"DD",x"7E",x"19",x"E6", -- 0x01F8
		x"07",x"C2",x"E8",x"2A",x"CD",x"38",x"4E",x"C3", -- 0x0200
		x"E8",x"2A",x"E5",x"21",x"D4",x"78",x"18",x"14", -- 0x0208
		x"DD",x"7E",x"01",x"E5",x"21",x"D4",x"78",x"E6", -- 0x0210
		x"C0",x"28",x"09",x"21",x"24",x"79",x"07",x"30", -- 0x0218
		x"03",x"21",x"54",x"79",x"C5",x"DD",x"4E",x"19", -- 0x0220
		x"06",x"00",x"09",x"C1",x"7E",x"E1",x"C9",x"E5", -- 0x0228
		x"21",x"24",x"79",x"18",x"EF",x"E5",x"21",x"54", -- 0x0230
		x"79",x"18",x"E9",x"3A",x"1C",x"E1",x"DD",x"77", -- 0x0238
		x"16",x"07",x"4F",x"06",x"00",x"21",x"AA",x"42", -- 0x0240
		x"09",x"7E",x"23",x"66",x"6F",x"56",x"23",x"3A", -- 0x0248
		x"03",x"E1",x"E6",x"1F",x"07",x"4F",x"09",x"C5", -- 0x0250
		x"3A",x"EF",x"E0",x"5E",x"06",x"EF",x"CB",x"57", -- 0x0258
		x"28",x"08",x"3E",x"10",x"93",x"D6",x"03",x"5F", -- 0x0260
		x"06",x"01",x"DD",x"70",x"0E",x"E6",x"03",x"83", -- 0x0268
		x"DD",x"77",x"14",x"DD",x"77",x"19",x"3A",x"0C", -- 0x0270
		x"E0",x"83",x"A2",x"23",x"86",x"DD",x"77",x"0F", -- 0x0278
		x"C1",x"21",x"73",x"43",x"09",x"7E",x"DD",x"77", -- 0x0280
		x"22",x"23",x"7E",x"DD",x"77",x"23",x"CD",x"26", -- 0x0288
		x"45",x"3A",x"EF",x"E0",x"E6",x"0F",x"C6",x"10", -- 0x0290
		x"DD",x"77",x"13",x"CD",x"10",x"42",x"DD",x"77", -- 0x0298
		x"0C",x"DD",x"34",x"03",x"C3",x"E8",x"2A",x"0C", -- 0x02A0
		x"0C",x"0E",x"B0",x"42",x"F1",x"42",x"32",x"43", -- 0x02A8
		x"7F",x"01",x"60",x"01",x"60",x"01",x"60",x"02", -- 0x02B0
		x"60",x"02",x"60",x"03",x"60",x"03",x"60",x"04", -- 0x02B8
		x"60",x"03",x"60",x"04",x"60",x"03",x"60",x"04", -- 0x02C0
		x"60",x"03",x"60",x"04",x"60",x"03",x"60",x"04", -- 0x02C8
		x"60",x"03",x"60",x"04",x"60",x"03",x"60",x"04", -- 0x02D0
		x"60",x"03",x"60",x"04",x"60",x"03",x"60",x"04", -- 0x02D8
		x"60",x"03",x"60",x"04",x"60",x"03",x"60",x"04", -- 0x02E0
		x"60",x"03",x"60",x"04",x"60",x"03",x"60",x"04", -- 0x02E8
		x"60",x"3F",x"01",x"60",x"01",x"60",x"01",x"60", -- 0x02F0
		x"01",x"60",x"01",x"60",x"01",x"60",x"01",x"60", -- 0x02F8
		x"01",x"60",x"01",x"60",x"02",x"60",x"03",x"60", -- 0x0300
		x"04",x"60",x"03",x"60",x"04",x"60",x"04",x"60", -- 0x0308
		x"04",x"60",x"04",x"60",x"04",x"60",x"04",x"60", -- 0x0310
		x"04",x"60",x"04",x"60",x"04",x"60",x"04",x"60", -- 0x0318
		x"04",x"60",x"04",x"60",x"04",x"60",x"04",x"60", -- 0x0320
		x"04",x"60",x"04",x"60",x"04",x"60",x"04",x"60", -- 0x0328
		x"04",x"60",x"3F",x"01",x"80",x"01",x"80",x"01", -- 0x0330
		x"80",x"01",x"80",x"01",x"80",x"01",x"80",x"01", -- 0x0338
		x"80",x"01",x"80",x"01",x"80",x"01",x"80",x"01", -- 0x0340
		x"80",x"01",x"80",x"01",x"80",x"01",x"80",x"01", -- 0x0348
		x"80",x"03",x"90",x"01",x"80",x"02",x"88",x"03", -- 0x0350
		x"90",x"04",x"9F",x"03",x"90",x"03",x"90",x"03", -- 0x0358
		x"90",x"04",x"9F",x"03",x"90",x"03",x"90",x"03", -- 0x0360
		x"90",x"04",x"9F",x"03",x"90",x"03",x"90",x"03", -- 0x0368
		x"90",x"04",x"9F",x"68",x"01",x"E0",x"01",x"1C", -- 0x0370
		x"02",x"58",x"02",x"E0",x"01",x"1C",x"02",x"1C", -- 0x0378
		x"02",x"58",x"02",x"1C",x"02",x"1C",x"02",x"58", -- 0x0380
		x"02",x"58",x"02",x"58",x"02",x"94",x"02",x"D0", -- 0x0388
		x"02",x"0C",x"03",x"1C",x"02",x"1C",x"02",x"58", -- 0x0390
		x"02",x"94",x"02",x"58",x"02",x"D0",x"02",x"48", -- 0x0398
		x"03",x"C0",x"03",x"D0",x"02",x"48",x"03",x"C0", -- 0x03A0
		x"03",x"B0",x"04",x"48",x"03",x"B0",x"04",x"80", -- 0x03A8
		x"07",x"80",x"07",x"CD",x"C5",x"43",x"DD",x"35", -- 0x03B0
		x"13",x"C2",x"E8",x"2A",x"DD",x"34",x"13",x"DD", -- 0x03B8
		x"34",x"03",x"C3",x"E8",x"2A",x"21",x"7D",x"46", -- 0x03C0
		x"DD",x"7E",x"14",x"CB",x"47",x"28",x"03",x"21", -- 0x03C8
		x"83",x"46",x"E6",x"0E",x"07",x"4F",x"06",x"00", -- 0x03D0
		x"DD",x"7E",x"16",x"07",x"5F",x"50",x"19",x"5E", -- 0x03D8
		x"23",x"56",x"EB",x"DD",x"34",x"15",x"DD",x"CB", -- 0x03E0
		x"15",x"46",x"28",x"02",x"CB",x"C9",x"06",x"00", -- 0x03E8
		x"09",x"4E",x"23",x"46",x"C3",x"FB",x"3A",x"CD", -- 0x03F0
		x"EC",x"50",x"CD",x"C5",x"43",x"DA",x"7D",x"44", -- 0x03F8
		x"DD",x"6E",x"22",x"DD",x"66",x"23",x"7D",x"B4", -- 0x0400
		x"CA",x"E8",x"2A",x"2B",x"DD",x"75",x"22",x"DD", -- 0x0408
		x"74",x"23",x"DD",x"35",x"13",x"C2",x"E8",x"2A", -- 0x0410
		x"DD",x"7E",x"16",x"4F",x"06",x"00",x"21",x"A7", -- 0x0418
		x"42",x"09",x"7E",x"DD",x"77",x"13",x"3A",x"C7", -- 0x0420
		x"E0",x"B7",x"C2",x"E8",x"2A",x"DD",x"CB",x"0D", -- 0x0428
		x"66",x"C2",x"E8",x"2A",x"DD",x"7E",x"19",x"E6", -- 0x0430
		x"0F",x"CD",x"F7",x"66",x"81",x"44",x"CA",x"45", -- 0x0438
		x"2E",x"45",x"FE",x"45",x"9C",x"44",x"D7",x"45", -- 0x0440
		x"4B",x"45",x"1B",x"46",x"B5",x"44",x"E4",x"45", -- 0x0448
		x"67",x"45",x"37",x"46",x"D7",x"44",x"F1",x"45", -- 0x0450
		x"84",x"45",x"4B",x"46",x"DD",x"72",x"21",x"7A", -- 0x0458
		x"FE",x"01",x"DD",x"7E",x"19",x"20",x"04",x"3C", -- 0x0460
		x"C3",x"6C",x"44",x"3D",x"E6",x"0F",x"DD",x"77", -- 0x0468
		x"19",x"DD",x"77",x"14",x"CD",x"10",x"42",x"DD", -- 0x0470
		x"77",x"0C",x"C3",x"E8",x"2A",x"CD",x"FD",x"64", -- 0x0478
		x"C9",x"CD",x"07",x"45",x"7D",x"11",x"66",x"46", -- 0x0480
		x"B7",x"C2",x"94",x"44",x"CB",x"49",x"CA",x"E8", -- 0x0488
		x"2A",x"C3",x"98",x"45",x"CB",x"49",x"C2",x"FF", -- 0x0490
		x"44",x"C3",x"CC",x"44",x"CD",x"07",x"45",x"11", -- 0x0498
		x"62",x"46",x"B7",x"20",x"08",x"CB",x"41",x"C2", -- 0x04A0
		x"E8",x"2A",x"C3",x"98",x"45",x"CB",x"41",x"CA", -- 0x04A8
		x"FF",x"44",x"C3",x"F7",x"44",x"CD",x"07",x"45", -- 0x04B0
		x"7D",x"11",x"5E",x"46",x"B7",x"20",x"08",x"CB", -- 0x04B8
		x"49",x"C2",x"E8",x"2A",x"C3",x"E8",x"44",x"CB", -- 0x04C0
		x"49",x"CA",x"FF",x"44",x"7C",x"0F",x"E6",x"F0", -- 0x04C8
		x"BD",x"D2",x"E8",x"2A",x"C3",x"FF",x"44",x"CD", -- 0x04D0
		x"07",x"45",x"11",x"6A",x"46",x"B7",x"20",x"12", -- 0x04D8
		x"CB",x"41",x"CA",x"E8",x"2A",x"C3",x"98",x"45", -- 0x04E0
		x"3A",x"0C",x"E0",x"07",x"E6",x"01",x"57",x"C3", -- 0x04E8
		x"5C",x"44",x"CB",x"41",x"C2",x"FF",x"44",x"7D", -- 0x04F0
		x"0F",x"E6",x"F0",x"BC",x"D2",x"E8",x"2A",x"EB", -- 0x04F8
		x"06",x"00",x"09",x"56",x"C3",x"5C",x"44",x"CD", -- 0x0500
		x"26",x"45",x"0E",x"00",x"7D",x"DD",x"96",x"0E", -- 0x0508
		x"30",x"03",x"0C",x"ED",x"44",x"E6",x"F0",x"6F", -- 0x0510
		x"7C",x"DD",x"96",x"0F",x"30",x"04",x"CB",x"C9", -- 0x0518
		x"ED",x"44",x"E6",x"F0",x"67",x"C9",x"2A",x"0E", -- 0x0520
		x"E1",x"7D",x"C6",x"08",x"6F",x"C9",x"CD",x"07", -- 0x0528
		x"45",x"BD",x"11",x"6F",x"46",x"79",x"C2",x"46", -- 0x0530
		x"45",x"FE",x"01",x"CA",x"E8",x"2A",x"FE",x"02", -- 0x0538
		x"CA",x"98",x"45",x"C3",x"BB",x"45",x"FE",x"01", -- 0x0540
		x"C3",x"9F",x"45",x"CD",x"07",x"45",x"BD",x"11", -- 0x0548
		x"60",x"46",x"79",x"C2",x"62",x"45",x"FE",x"03", -- 0x0550
		x"CA",x"E8",x"2A",x"B7",x"CA",x"98",x"45",x"C3", -- 0x0558
		x"BB",x"45",x"FE",x"03",x"C3",x"9F",x"45",x"CD", -- 0x0560
		x"07",x"45",x"BD",x"11",x"75",x"46",x"79",x"C2", -- 0x0568
		x"7F",x"45",x"FE",x"02",x"CA",x"E8",x"2A",x"FE", -- 0x0570
		x"01",x"CA",x"98",x"45",x"C3",x"BB",x"45",x"FE", -- 0x0578
		x"02",x"C3",x"9F",x"45",x"CD",x"07",x"45",x"BD", -- 0x0580
		x"11",x"68",x"46",x"79",x"C2",x"9E",x"45",x"B7", -- 0x0588
		x"CA",x"E8",x"2A",x"FE",x"03",x"C2",x"BB",x"45", -- 0x0590
		x"DD",x"56",x"21",x"C3",x"5C",x"44",x"B7",x"C2", -- 0x0598
		x"BB",x"45",x"7D",x"0F",x"E6",x"F0",x"BC",x"CA", -- 0x05A0
		x"E8",x"2A",x"30",x"0E",x"7C",x"0F",x"E6",x"F0", -- 0x05A8
		x"67",x"BD",x"DA",x"E8",x"2A",x"CA",x"E8",x"2A", -- 0x05B0
		x"18",x"01",x"6F",x"EB",x"CB",x"01",x"06",x"00", -- 0x05B8
		x"09",x"7A",x"BB",x"38",x"01",x"23",x"56",x"C3", -- 0x05C0
		x"5C",x"44",x"CD",x"07",x"45",x"79",x"EE",x"01", -- 0x05C8
		x"4F",x"11",x"60",x"46",x"C3",x"51",x"46",x"CD", -- 0x05D0
		x"07",x"45",x"79",x"EE",x"01",x"4F",x"11",x"6F", -- 0x05D8
		x"46",x"C3",x"3D",x"46",x"CD",x"07",x"45",x"79", -- 0x05E0
		x"EE",x"01",x"4F",x"11",x"68",x"46",x"C3",x"21", -- 0x05E8
		x"46",x"CD",x"07",x"45",x"79",x"EE",x"01",x"4F", -- 0x05F0
		x"11",x"75",x"46",x"C3",x"04",x"46",x"CD",x"07", -- 0x05F8
		x"45",x"11",x"6F",x"46",x"79",x"FE",x"02",x"28", -- 0x0600
		x"0C",x"FE",x"01",x"20",x"0B",x"7D",x"BC",x"D2", -- 0x0608
		x"E8",x"2A",x"C3",x"BB",x"45",x"C3",x"98",x"45", -- 0x0610
		x"C3",x"BB",x"45",x"CD",x"07",x"45",x"11",x"60", -- 0x0618
		x"46",x"79",x"B7",x"28",x"0C",x"FE",x"03",x"20", -- 0x0620
		x"0B",x"7C",x"BD",x"D2",x"E8",x"2A",x"C3",x"BB", -- 0x0628
		x"45",x"C3",x"98",x"45",x"C3",x"BB",x"45",x"CD", -- 0x0630
		x"07",x"45",x"11",x"75",x"46",x"79",x"FE",x"01", -- 0x0638
		x"CA",x"15",x"46",x"FE",x"02",x"C2",x"18",x"46", -- 0x0640
		x"C3",x"0D",x"46",x"CD",x"07",x"45",x"11",x"68", -- 0x0648
		x"46",x"79",x"FE",x"03",x"CA",x"31",x"46",x"B7", -- 0x0650
		x"C2",x"34",x"46",x"C3",x"29",x"46",x"01",x"02", -- 0x0658
		x"01",x"02",x"02",x"02",x"01",x"01",x"02",x"01", -- 0x0660
		x"02",x"01",x"01",x"01",x"02",x"02",x"01",x"02", -- 0x0668
		x"02",x"01",x"02",x"02",x"01",x"01",x"01",x"02", -- 0x0670
		x"01",x"01",x"02",x"02",x"02",x"89",x"46",x"C9", -- 0x0678
		x"46",x"09",x"47",x"A9",x"46",x"E9",x"46",x"29", -- 0x0680
		x"47",x"01",x"00",x"01",x"00",x"01",x"FF",x"01", -- 0x0688
		x"FF",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x0690
		x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"01",x"FF", -- 0x0698
		x"01",x"00",x"01",x"00",x"01",x"01",x"01",x"01", -- 0x06A0
		x"01",x"01",x"00",x"01",x"FF",x"00",x"FF",x"01", -- 0x06A8
		x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x06B0
		x"FF",x"FF",x"00",x"FF",x"01",x"00",x"01",x"FF", -- 0x06B8
		x"01",x"00",x"01",x"01",x"01",x"01",x"00",x"01", -- 0x06C0
		x"01",x"02",x"00",x"01",x"00",x"02",x"FE",x"01", -- 0x06C8
		x"FF",x"00",x"FE",x"00",x"FF",x"FE",x"FE",x"FF", -- 0x06D0
		x"FF",x"FE",x"00",x"FF",x"00",x"FE",x"02",x"FF", -- 0x06D8
		x"01",x"00",x"02",x"00",x"01",x"02",x"02",x"01", -- 0x06E0
		x"01",x"01",x"00",x"02",x"FF",x"00",x"FF",x"01", -- 0x06E8
		x"FE",x"00",x"FF",x"FF",x"FE",x"FF",x"00",x"FE", -- 0x06F0
		x"FF",x"FF",x"00",x"FE",x"01",x"00",x"01",x"FF", -- 0x06F8
		x"02",x"00",x"01",x"01",x"02",x"01",x"00",x"02", -- 0x0700
		x"01",x"02",x"00",x"02",x"00",x"02",x"FE",x"02", -- 0x0708
		x"FE",x"00",x"FE",x"00",x"FE",x"FE",x"FE",x"FE", -- 0x0710
		x"FE",x"FE",x"00",x"FE",x"00",x"FE",x"02",x"FE", -- 0x0718
		x"02",x"00",x"02",x"00",x"02",x"02",x"02",x"02", -- 0x0720
		x"02",x"02",x"FF",x"02",x"FF",x"01",x"FE",x"01", -- 0x0728
		x"FE",x"FF",x"FE",x"FF",x"FE",x"FE",x"FF",x"FE", -- 0x0730
		x"FF",x"FE",x"01",x"FE",x"01",x"FF",x"02",x"FF", -- 0x0738
		x"02",x"01",x"02",x"01",x"02",x"02",x"01",x"02", -- 0x0740
		x"01",x"CD",x"82",x"36",x"DD",x"CB",x"1A",x"46", -- 0x0748
		x"C2",x"BD",x"47",x"DD",x"36",x"19",x"00",x"DD", -- 0x0750
		x"36",x"0C",x"68",x"01",x"1F",x"80",x"CD",x"E5", -- 0x0758
		x"47",x"3A",x"0C",x"E0",x"6F",x"3A",x"F0",x"E0", -- 0x0760
		x"85",x"32",x"F0",x"E0",x"CB",x"57",x"CA",x"96", -- 0x0768
		x"47",x"DD",x"36",x"0E",x"EF",x"DD",x"36",x"02", -- 0x0770
		x"03",x"21",x"8E",x"91",x"DD",x"75",x"10",x"DD", -- 0x0778
		x"74",x"11",x"7E",x"DD",x"77",x"14",x"DD",x"7E", -- 0x0780
		x"1A",x"0F",x"E6",x"80",x"DD",x"B6",x"02",x"DD", -- 0x0788
		x"77",x"02",x"DD",x"34",x"03",x"C9",x"DD",x"36", -- 0x0790
		x"0E",x"01",x"DD",x"36",x"02",x"0B",x"18",x"D9", -- 0x0798
		x"DD",x"36",x"19",x"0C",x"DD",x"36",x"0C",x"64", -- 0x07A0
		x"DD",x"36",x"0E",x"01",x"DD",x"36",x"02",x"80", -- 0x07A8
		x"DD",x"36",x"16",x"40",x"DD",x"36",x"09",x"02", -- 0x07B0
		x"21",x"DE",x"90",x"18",x"BF",x"01",x"1F",x"08", -- 0x07B8
		x"CD",x"E5",x"47",x"3A",x"0C",x"E0",x"6F",x"3A", -- 0x07C0
		x"F0",x"E0",x"85",x"32",x"F0",x"E0",x"CB",x"57", -- 0x07C8
		x"CA",x"A0",x"47",x"DD",x"36",x"19",x"04",x"DD", -- 0x07D0
		x"36",x"0C",x"6C",x"DD",x"36",x"0E",x"EF",x"DD", -- 0x07D8
		x"36",x"02",x"89",x"18",x"CB",x"CD",x"D4",x"56", -- 0x07E0
		x"A1",x"80",x"DD",x"77",x"0F",x"C9",x"DD",x"7E", -- 0x07E8
		x"02",x"CB",x"7F",x"C2",x"FF",x"47",x"CD",x"9A", -- 0x07F0
		x"4A",x"D2",x"59",x"3C",x"C3",x"9E",x"48",x"DD", -- 0x07F8
		x"6E",x"10",x"DD",x"66",x"11",x"23",x"CB",x"5F", -- 0x0800
		x"7E",x"C4",x"90",x"39",x"47",x"DD",x"86",x"0E", -- 0x0808
		x"DD",x"77",x"0E",x"3A",x"C7",x"E0",x"B7",x"CA", -- 0x0810
		x"24",x"48",x"78",x"DD",x"86",x"0E",x"DD",x"77", -- 0x0818
		x"0E",x"C3",x"59",x"3C",x"DD",x"35",x"14",x"C2", -- 0x0820
		x"59",x"3C",x"23",x"7E",x"B7",x"28",x"0C",x"DD", -- 0x0828
		x"77",x"14",x"DD",x"75",x"10",x"DD",x"74",x"11", -- 0x0830
		x"C3",x"59",x"3C",x"21",x"45",x"91",x"DD",x"75", -- 0x0838
		x"10",x"DD",x"74",x"11",x"7E",x"DD",x"77",x"14", -- 0x0840
		x"DD",x"34",x"03",x"C3",x"59",x"3C",x"CD",x"9A", -- 0x0848
		x"4A",x"D2",x"59",x"3C",x"3A",x"0C",x"E0",x"E6", -- 0x0850
		x"07",x"3C",x"DD",x"77",x"14",x"DD",x"34",x"03", -- 0x0858
		x"C3",x"59",x"3C",x"DD",x"7E",x"09",x"DD",x"86", -- 0x0860
		x"0F",x"DD",x"77",x"0F",x"FE",x"80",x"DA",x"E8", -- 0x0868
		x"2A",x"DD",x"35",x"14",x"C2",x"E8",x"2A",x"3A", -- 0x0870
		x"C7",x"E0",x"B7",x"C2",x"59",x"3C",x"21",x"8E", -- 0x0878
		x"91",x"DD",x"75",x"10",x"DD",x"74",x"11",x"7E", -- 0x0880
		x"DD",x"77",x"14",x"DD",x"34",x"03",x"C3",x"E8", -- 0x0888
		x"2A",x"CD",x"9A",x"4A",x"D2",x"59",x"3C",x"3A", -- 0x0890
		x"0F",x"E1",x"FE",x"70",x"30",x"4E",x"21",x"94", -- 0x0898
		x"92",x"3A",x"0E",x"E1",x"DD",x"CB",x"02",x"5E", -- 0x08A0
		x"20",x"0A",x"DD",x"96",x"0E",x"D2",x"D5",x"48", -- 0x08A8
		x"ED",x"44",x"18",x"06",x"DD",x"96",x"0E",x"DA", -- 0x08B0
		x"D5",x"48",x"E6",x"F0",x"FE",x"B0",x"DA",x"D5", -- 0x08B8
		x"48",x"21",x"2C",x"9B",x"FE",x"E0",x"D2",x"D5", -- 0x08C0
		x"48",x"0F",x"4F",x"06",x"00",x"21",x"15",x"92", -- 0x08C8
		x"09",x"7E",x"23",x"66",x"6F",x"DD",x"75",x"10", -- 0x08D0
		x"DD",x"74",x"11",x"7E",x"DD",x"77",x"14",x"CD", -- 0x08D8
		x"35",x"42",x"DD",x"77",x"0C",x"DD",x"36",x"03", -- 0x08E0
		x"09",x"C3",x"59",x"3C",x"DD",x"34",x"03",x"21", -- 0x08E8
		x"5C",x"96",x"DD",x"75",x"10",x"DD",x"74",x"11", -- 0x08F0
		x"7E",x"DD",x"77",x"14",x"DD",x"36",x"13",x"02", -- 0x08F8
		x"C3",x"59",x"3C",x"CD",x"EC",x"50",x"CD",x"9A", -- 0x0900
		x"4A",x"D2",x"59",x"3C",x"DD",x"35",x"13",x"28", -- 0x0908
		x"10",x"21",x"B9",x"96",x"DD",x"75",x"10",x"DD", -- 0x0910
		x"74",x"11",x"7E",x"DD",x"77",x"14",x"C3",x"59", -- 0x0918
		x"3C",x"DD",x"34",x"03",x"3A",x"0F",x"E1",x"FE", -- 0x0920
		x"70",x"38",x"5C",x"3A",x"0E",x"E1",x"DD",x"CB", -- 0x0928
		x"02",x"5E",x"20",x"07",x"DD",x"96",x"0E",x"38", -- 0x0930
		x"4E",x"18",x"07",x"DD",x"96",x"0E",x"30",x"47", -- 0x0938
		x"ED",x"44",x"E6",x"F0",x"47",x"3A",x"0F",x"E1", -- 0x0940
		x"DD",x"96",x"0F",x"DC",x"90",x"39",x"E6",x"F0", -- 0x0948
		x"B8",x"30",x"01",x"78",x"21",x"1A",x"9E",x"FE", -- 0x0950
		x"E0",x"30",x"15",x"21",x"16",x"93",x"FE",x"90", -- 0x0958
		x"38",x"0E",x"D6",x"90",x"0F",x"4F",x"06",x"00", -- 0x0960
		x"21",x"21",x"92",x"09",x"7E",x"23",x"66",x"6F", -- 0x0968
		x"DD",x"75",x"10",x"DD",x"74",x"11",x"23",x"7E", -- 0x0970
		x"DD",x"77",x"14",x"CD",x"35",x"42",x"DD",x"77", -- 0x0978
		x"0C",x"DD",x"34",x"03",x"C3",x"59",x"3C",x"21", -- 0x0980
		x"1A",x"9E",x"DD",x"75",x"10",x"DD",x"74",x"11", -- 0x0988
		x"7E",x"DD",x"77",x"14",x"DD",x"36",x"13",x"02", -- 0x0990
		x"C3",x"59",x"3C",x"CD",x"9A",x"4A",x"D2",x"59", -- 0x0998
		x"3C",x"DD",x"35",x"13",x"28",x"10",x"21",x"7F", -- 0x09A0
		x"9C",x"DD",x"75",x"10",x"DD",x"74",x"11",x"7E", -- 0x09A8
		x"DD",x"77",x"14",x"C3",x"59",x"3C",x"DD",x"36", -- 0x09B0
		x"14",x"FF",x"C3",x"59",x"3C",x"CD",x"EC",x"50", -- 0x09B8
		x"CD",x"9A",x"4A",x"D2",x"59",x"3C",x"21",x"7B", -- 0x09C0
		x"9F",x"3A",x"0E",x"E1",x"DD",x"CB",x"02",x"5E", -- 0x09C8
		x"20",x"0A",x"DD",x"96",x"0E",x"D2",x"E2",x"49", -- 0x09D0
		x"ED",x"44",x"18",x"0C",x"DD",x"96",x"0E",x"D2", -- 0x09D8
		x"E8",x"49",x"CD",x"1F",x"4B",x"C3",x"EB",x"49", -- 0x09E0
		x"CD",x"EB",x"4A",x"DD",x"7E",x"19",x"E6",x"0C", -- 0x09E8
		x"07",x"C6",x"10",x"DD",x"77",x"19",x"DD",x"36", -- 0x09F0
		x"16",x"01",x"DD",x"34",x"03",x"C3",x"59",x"3C", -- 0x09F8
		x"CD",x"EC",x"50",x"CD",x"E3",x"4A",x"D2",x"0D", -- 0x0A00
		x"4A",x"DD",x"36",x"14",x"FF",x"DD",x"35",x"16", -- 0x0A08
		x"C2",x"59",x"3C",x"DD",x"36",x"16",x"02",x"DD", -- 0x0A10
		x"7E",x"19",x"4F",x"DD",x"CB",x"02",x"5E",x"20", -- 0x0A18
		x"0F",x"E6",x"07",x"20",x"08",x"79",x"E6",x"38", -- 0x0A20
		x"F6",x"07",x"4F",x"18",x"0F",x"0D",x"18",x"0C", -- 0x0A28
		x"3C",x"E6",x"07",x"20",x"06",x"79",x"E6",x"38", -- 0x0A30
		x"4F",x"18",x"01",x"0C",x"DD",x"71",x"19",x"CD", -- 0x0A38
		x"35",x"42",x"DD",x"77",x"0C",x"C3",x"59",x"3C", -- 0x0A40
		x"CD",x"EC",x"50",x"CD",x"9A",x"4A",x"D2",x"59", -- 0x0A48
		x"3C",x"21",x"E9",x"9E",x"3A",x"0F",x"E1",x"DD", -- 0x0A50
		x"BE",x"0F",x"D2",x"E2",x"49",x"21",x"7B",x"9F", -- 0x0A58
		x"3A",x"0E",x"E1",x"DD",x"CB",x"02",x"5E",x"20", -- 0x0A60
		x"09",x"DD",x"96",x"0E",x"DA",x"E2",x"49",x"C3", -- 0x0A68
		x"E8",x"49",x"DD",x"96",x"0E",x"D2",x"E2",x"49", -- 0x0A70
		x"ED",x"44",x"C3",x"E8",x"49",x"CD",x"EC",x"50", -- 0x0A78
		x"DD",x"6E",x"10",x"DD",x"66",x"11",x"23",x"7E", -- 0x0A80
		x"ED",x"44",x"4F",x"23",x"7E",x"DD",x"CB",x"02", -- 0x0A88
		x"5E",x"CC",x"90",x"39",x"CD",x"C0",x"4A",x"C3", -- 0x0A90
		x"06",x"4A",x"DD",x"6E",x"10",x"DD",x"66",x"11", -- 0x0A98
		x"23",x"7E",x"DD",x"CB",x"02",x"5E",x"28",x"04", -- 0x0AA0
		x"ED",x"44",x"E6",x"0F",x"DD",x"77",x"19",x"CD", -- 0x0AA8
		x"10",x"42",x"DD",x"77",x"0C",x"23",x"4E",x"23", -- 0x0AB0
		x"7E",x"DD",x"CB",x"02",x"5E",x"C4",x"90",x"39", -- 0x0AB8
		x"47",x"E5",x"CD",x"E4",x"3C",x"E1",x"DD",x"35", -- 0x0AC0
		x"14",x"C2",x"DA",x"4A",x"23",x"7E",x"B7",x"28", -- 0x0AC8
		x"0B",x"DD",x"77",x"14",x"DD",x"75",x"10",x"DD", -- 0x0AD0
		x"74",x"11",x"B7",x"C9",x"3A",x"C7",x"E0",x"B7", -- 0x0AD8
		x"C0",x"37",x"C9",x"DD",x"6E",x"10",x"DD",x"66", -- 0x0AE0
		x"11",x"18",x"CA",x"E6",x"F0",x"FE",x"70",x"38", -- 0x0AE8
		x"02",x"3E",x"70",x"0F",x"4F",x"06",x"00",x"21", -- 0x0AF0
		x"A3",x"9E",x"09",x"3A",x"0F",x"E1",x"DD",x"96", -- 0x0AF8
		x"0F",x"DC",x"90",x"39",x"E6",x"F0",x"0F",x"0F", -- 0x0B00
		x"0F",x"0F",x"FE",x"08",x"38",x"04",x"0E",x"04", -- 0x0B08
		x"18",x"05",x"4F",x"09",x"7E",x"07",x"4F",x"21", -- 0x0B10
		x"E3",x"9E",x"09",x"7E",x"23",x"66",x"6F",x"DD", -- 0x0B18
		x"75",x"10",x"DD",x"74",x"11",x"7E",x"DD",x"77", -- 0x0B20
		x"14",x"C9",x"DD",x"CB",x"01",x"66",x"CA",x"38", -- 0x0B28
		x"4B",x"DD",x"CB",x"01",x"56",x"CA",x"55",x"4D", -- 0x0B30
		x"CD",x"EC",x"50",x"DD",x"CB",x"01",x"5E",x"C2", -- 0x0B38
		x"F2",x"40",x"DD",x"CB",x"02",x"56",x"C2",x"CE", -- 0x0B40
		x"4D",x"DD",x"7E",x"19",x"B7",x"CA",x"C0",x"4C", -- 0x0B48
		x"FE",x"08",x"CA",x"9E",x"4B",x"0E",x"04",x"DD", -- 0x0B50
		x"CB",x"02",x"5E",x"28",x"02",x"0E",x"0C",x"B9", -- 0x0B58
		x"C2",x"E3",x"4C",x"3A",x"C7",x"E0",x"B7",x"21", -- 0x0B60
		x"DE",x"87",x"3E",x"0F",x"C2",x"57",x"4C",x"21", -- 0x0B68
		x"BE",x"87",x"79",x"FE",x"04",x"20",x"07",x"DD", -- 0x0B70
		x"7E",x"0E",x"D6",x"10",x"18",x"05",x"3E",x"E0", -- 0x0B78
		x"DD",x"96",x"0E",x"DA",x"50",x"4C",x"0F",x"0F", -- 0x0B80
		x"0F",x"0F",x"E6",x"0F",x"FE",x"08",x"DA",x"50", -- 0x0B88
		x"4C",x"21",x"DE",x"87",x"FE",x"0F",x"D2",x"57", -- 0x0B90
		x"4C",x"D6",x"07",x"C3",x"40",x"4C",x"DD",x"34", -- 0x0B98
		x"13",x"0E",x"00",x"DD",x"CB",x"0D",x"66",x"3A", -- 0x0BA0
		x"0F",x"E1",x"20",x"0A",x"DD",x"96",x"0F",x"30", -- 0x0BA8
		x"0C",x"0C",x"ED",x"44",x"18",x"07",x"5F",x"DD", -- 0x0BB0
		x"7E",x"0F",x"ED",x"44",x"83",x"5F",x"3A",x"0E", -- 0x0BB8
		x"E1",x"C6",x"08",x"DD",x"96",x"0E",x"30",x"04", -- 0x0BC0
		x"ED",x"44",x"CB",x"C9",x"57",x"21",x"3E",x"7C", -- 0x0BC8
		x"DD",x"CB",x"02",x"5E",x"28",x"03",x"21",x"42", -- 0x0BD0
		x"7C",x"DD",x"7E",x"02",x"E6",x"03",x"06",x"00", -- 0x0BD8
		x"09",x"BE",x"21",x"BE",x"87",x"20",x"69",x"21", -- 0x0BE0
		x"DE",x"87",x"7B",x"DD",x"CB",x"01",x"56",x"20", -- 0x0BE8
		x"5F",x"7A",x"0F",x"0F",x"0F",x"0F",x"E6",x"0F", -- 0x0BF0
		x"57",x"7B",x"0F",x"0F",x"0F",x"0F",x"E6",x"0F", -- 0x0BF8
		x"5F",x"21",x"BE",x"87",x"FE",x"07",x"38",x"48", -- 0x0C00
		x"21",x"DE",x"87",x"FE",x"0F",x"30",x"48",x"7A", -- 0x0C08
		x"BB",x"30",x"02",x"53",x"5F",x"4A",x"7A",x"CB", -- 0x0C10
		x"3F",x"BB",x"30",x"04",x"47",x"7B",x"90",x"5F", -- 0x0C18
		x"79",x"FE",x"06",x"21",x"BE",x"87",x"38",x"28", -- 0x0C20
		x"21",x"DE",x"87",x"D6",x"06",x"FE",x"09",x"30", -- 0x0C28
		x"26",x"07",x"4F",x"06",x"00",x"21",x"E9",x"4C", -- 0x0C30
		x"09",x"7E",x"23",x"66",x"6F",x"50",x"19",x"7E", -- 0x0C38
		x"DD",x"77",x"20",x"21",x"A8",x"87",x"CD",x"09", -- 0x0C40
		x"41",x"7E",x"23",x"66",x"6F",x"C3",x"5C",x"4C", -- 0x0C48
		x"AF",x"DD",x"77",x"20",x"C3",x"5C",x"4C",x"3E", -- 0x0C50
		x"08",x"DD",x"77",x"20",x"DD",x"7E",x"02",x"E6", -- 0x0C58
		x"03",x"E2",x"66",x"4C",x"EE",x"03",x"DD",x"CB", -- 0x0C60
		x"02",x"5E",x"28",x"09",x"DD",x"CB",x"02",x"4E", -- 0x0C68
		x"C2",x"75",x"4C",x"EE",x"02",x"FE",x"02",x"38", -- 0x0C70
		x"02",x"D6",x"02",x"CD",x"09",x"41",x"7E",x"23", -- 0x0C78
		x"66",x"6F",x"AF",x"DD",x"77",x"15",x"7E",x"DD", -- 0x0C80
		x"77",x"16",x"23",x"CD",x"63",x"40",x"CD",x"2F", -- 0x0C88
		x"42",x"DD",x"77",x"0C",x"23",x"DD",x"75",x"1E", -- 0x0C90
		x"DD",x"74",x"1F",x"DD",x"CB",x"02",x"D6",x"DD", -- 0x0C98
		x"56",x"19",x"DD",x"5E",x"01",x"7A",x"E6",x"03", -- 0x0CA0
		x"28",x"04",x"CB",x"CB",x"18",x"08",x"CB",x"8B", -- 0x0CA8
		x"CB",x"43",x"20",x"05",x"CB",x"C3",x"DD",x"73", -- 0x0CB0
		x"01",x"CD",x"3A",x"40",x"D8",x"C3",x"E8",x"2A", -- 0x0CB8
		x"3A",x"C7",x"E0",x"B7",x"20",x"08",x"DD",x"7E", -- 0x0CC0
		x"0F",x"FE",x"80",x"D2",x"D7",x"4C",x"01",x"02", -- 0x0CC8
		x"00",x"CD",x"F8",x"3C",x"C3",x"59",x"3C",x"CD", -- 0x0CD0
		x"38",x"4E",x"21",x"BE",x"87",x"D2",x"57",x"4C", -- 0x0CD8
		x"C3",x"A1",x"4B",x"DD",x"7E",x"20",x"C3",x"43", -- 0x0CE0
		x"4C",x"FB",x"4C",x"01",x"4D",x"08",x"4D",x"10", -- 0x0CE8
		x"4D",x"19",x"4D",x"23",x"4D",x"2E",x"4D",x"3A", -- 0x0CF0
		x"4D",x"47",x"4D",x"00",x"00",x"00",x"00",x"00", -- 0x0CF8
		x"01",x"00",x"00",x"00",x"00",x"01",x"01",x"02", -- 0x0D00
		x"01",x"01",x"01",x"01",x"02",x"02",x"03",x"03", -- 0x0D08
		x"02",x"02",x"02",x"02",x"03",x"03",x"03",x"04", -- 0x0D10
		x"05",x"03",x"03",x"03",x"03",x"04",x"04",x"04", -- 0x0D18
		x"05",x"05",x"06",x"04",x"04",x"04",x"04",x"05", -- 0x0D20
		x"05",x"05",x"06",x"06",x"07",x"07",x"05",x"05", -- 0x0D28
		x"05",x"05",x"05",x"06",x"06",x"07",x"07",x"08", -- 0x0D30
		x"08",x"08",x"06",x"06",x"06",x"06",x"06",x"07", -- 0x0D38
		x"07",x"07",x"08",x"08",x"08",x"08",x"08",x"07", -- 0x0D40
		x"07",x"07",x"07",x"07",x"08",x"08",x"08",x"08", -- 0x0D48
		x"08",x"08",x"08",x"08",x"08",x"DD",x"7E",x"19", -- 0x0D50
		x"FE",x"10",x"30",x"0C",x"E6",x"0C",x"07",x"C6", -- 0x0D58
		x"10",x"4F",x"DD",x"36",x"16",x"04",x"18",x"2B", -- 0x0D60
		x"4F",x"DD",x"35",x"16",x"C2",x"A0",x"4D",x"DD", -- 0x0D68
		x"36",x"16",x"04",x"DD",x"CB",x"02",x"5E",x"20", -- 0x0D70
		x"09",x"3C",x"E6",x"07",x"28",x"09",x"0C",x"C3", -- 0x0D78
		x"93",x"4D",x"3D",x"E6",x"07",x"20",x"0B",x"DD", -- 0x0D80
		x"CB",x"02",x"E6",x"79",x"E6",x"38",x"0F",x"4F", -- 0x0D88
		x"18",x"01",x"0D",x"DD",x"71",x"19",x"CD",x"2F", -- 0x0D90
		x"42",x"DD",x"77",x"0C",x"DD",x"CB",x"01",x"9E", -- 0x0D98
		x"01",x"02",x"00",x"DD",x"CB",x"02",x"5E",x"28", -- 0x0DA0
		x"03",x"01",x"FE",x"FF",x"DD",x"CB",x"0D",x"66", -- 0x0DA8
		x"C2",x"CB",x"66",x"CB",x"79",x"DD",x"7E",x"0E", -- 0x0DB0
		x"20",x"0A",x"81",x"DD",x"77",x"0E",x"DA",x"CB", -- 0x0DB8
		x"66",x"C3",x"E8",x"2A",x"81",x"DD",x"77",x"0E", -- 0x0DC0
		x"D2",x"CB",x"66",x"C3",x"E8",x"2A",x"DD",x"6E", -- 0x0DC8
		x"1E",x"DD",x"66",x"1F",x"E5",x"CD",x"3A",x"40", -- 0x0DD0
		x"E1",x"D8",x"23",x"23",x"3A",x"C7",x"E0",x"B7", -- 0x0DD8
		x"C2",x"E8",x"2A",x"DD",x"35",x"16",x"C2",x"E8", -- 0x0DE0
		x"2A",x"7E",x"B7",x"CA",x"0D",x"4E",x"DD",x"77", -- 0x0DE8
		x"16",x"23",x"CD",x"63",x"40",x"E6",x"03",x"28", -- 0x0DF0
		x"04",x"DD",x"CB",x"01",x"CE",x"CD",x"10",x"42", -- 0x0DF8
		x"DD",x"77",x"0C",x"23",x"DD",x"75",x"1E",x"DD", -- 0x0E00
		x"74",x"1F",x"C3",x"E8",x"2A",x"DD",x"7E",x"19", -- 0x0E08
		x"5F",x"FE",x"08",x"20",x"08",x"DD",x"CB",x"01", -- 0x0E10
		x"86",x"DD",x"CB",x"01",x"D6",x"7B",x"E6",x"0C", -- 0x0E18
		x"E2",x"25",x"4E",x"EE",x"0C",x"0F",x"0F",x"5F", -- 0x0E20
		x"DD",x"7E",x"02",x"E6",x"F8",x"B3",x"DD",x"77", -- 0x0E28
		x"02",x"DD",x"CB",x"01",x"8E",x"C3",x"E8",x"2A", -- 0x0E30
		x"DD",x"6E",x"10",x"DD",x"66",x"11",x"7E",x"FE", -- 0x0E38
		x"FF",x"C8",x"DD",x"77",x"12",x"3A",x"C7",x"E0", -- 0x0E40
		x"B7",x"C0",x"23",x"DD",x"75",x"10",x"DD",x"74", -- 0x0E48
		x"11",x"DD",x"36",x"03",x"01",x"01",x"68",x"4E", -- 0x0E50
		x"C5",x"CD",x"F7",x"66",x"24",x"39",x"B2",x"3B", -- 0x0E58
		x"A9",x"3B",x"06",x"3F",x"2D",x"3F",x"72",x"41", -- 0x0E60
		x"37",x"C9",x"DD",x"7E",x"14",x"B7",x"28",x"04", -- 0x0E68
		x"DD",x"35",x"14",x"C9",x"DD",x"36",x"18",x"01", -- 0x0E70
		x"AF",x"DD",x"77",x"13",x"DD",x"77",x"0A",x"DD", -- 0x0E78
		x"77",x"24",x"DD",x"77",x"25",x"DD",x"7E",x"08", -- 0x0E80
		x"57",x"CB",x"7F",x"01",x"A2",x"08",x"28",x"0F", -- 0x0E88
		x"E6",x"18",x"0F",x"0F",x"0F",x"4F",x"06",x"00", -- 0x0E90
		x"21",x"CA",x"4E",x"09",x"4E",x"06",x"00",x"DD", -- 0x0E98
		x"71",x"0C",x"79",x"D6",x"02",x"DD",x"77",x"2C", -- 0x0EA0
		x"DD",x"70",x"19",x"CD",x"82",x"36",x"3A",x"0C", -- 0x0EA8
		x"E0",x"07",x"07",x"E6",x"1F",x"C6",x"10",x"DD", -- 0x0EB0
		x"77",x"04",x"DD",x"34",x"03",x"DD",x"7E",x"08", -- 0x0EB8
		x"07",x"E6",x"01",x"CD",x"F7",x"66",x"CD",x"4E", -- 0x0EC0
		x"D9",x"4E",x"3E",x"3A",x"82",x"21",x"C2",x"B1", -- 0x0EC8
		x"CD",x"0B",x"50",x"DD",x"36",x"17",x"30",x"18", -- 0x0ED0
		x"0F",x"DD",x"7E",x"02",x"E6",x"07",x"FE",x"05", -- 0x0ED8
		x"20",x"06",x"CD",x"01",x"4F",x"DD",x"77",x"0E", -- 0x0EE0
		x"DD",x"7E",x"0E",x"DD",x"77",x"2E",x"DD",x"7E", -- 0x0EE8
		x"0F",x"C6",x"10",x"DD",x"77",x"2F",x"DD",x"7E", -- 0x0EF0
		x"0D",x"30",x"02",x"EE",x"10",x"DD",x"77",x"2D", -- 0x0EF8
		x"C9",x"3A",x"F1",x"E0",x"3C",x"32",x"F1",x"E0", -- 0x0F00
		x"0F",x"06",x"18",x"30",x"02",x"06",x"48",x"2A", -- 0x0F08
		x"EF",x"E0",x"3A",x"0C",x"E0",x"84",x"85",x"07", -- 0x0F10
		x"07",x"2F",x"22",x"EF",x"E0",x"21",x"E0",x"E0", -- 0x0F18
		x"34",x"86",x"E6",x"7F",x"80",x"C9",x"DD",x"7E", -- 0x0F20
		x"08",x"07",x"E6",x"01",x"CD",x"F7",x"66",x"33", -- 0x0F28
		x"4F",x"B0",x"4F",x"CD",x"EC",x"50",x"DD",x"7E", -- 0x0F30
		x"13",x"B7",x"28",x"0B",x"3D",x"CA",x"81",x"4F", -- 0x0F38
		x"3D",x"28",x"04",x"3D",x"CA",x"81",x"4F",x"3A", -- 0x0F40
		x"C7",x"E0",x"21",x"40",x"01",x"B7",x"20",x"03", -- 0x0F48
		x"21",x"80",x"01",x"CD",x"7A",x"50",x"3A",x"C7", -- 0x0F50
		x"E0",x"B7",x"C2",x"D2",x"4F",x"DD",x"35",x"17", -- 0x0F58
		x"C2",x"D2",x"4F",x"DD",x"CB",x"01",x"E6",x"DD", -- 0x0F60
		x"7E",x"13",x"B7",x"28",x"04",x"FE",x"02",x"20", -- 0x0F68
		x"09",x"DD",x"34",x"13",x"CD",x"08",x"50",x"C3", -- 0x0F70
		x"D2",x"4F",x"DD",x"36",x"17",x"FF",x"C3",x"D2", -- 0x0F78
		x"4F",x"CD",x"35",x"50",x"DD",x"35",x"16",x"C2", -- 0x0F80
		x"D2",x"4F",x"DD",x"6E",x"10",x"DD",x"66",x"11", -- 0x0F88
		x"23",x"23",x"7E",x"B7",x"28",x"06",x"CD",x"0C", -- 0x0F90
		x"50",x"C3",x"D2",x"4F",x"DD",x"7E",x"13",x"FE", -- 0x0F98
		x"01",x"06",x"50",x"28",x"02",x"06",x"FF",x"DD", -- 0x0FA0
		x"70",x"17",x"DD",x"34",x"13",x"C3",x"D2",x"4F", -- 0x0FA8
		x"CD",x"D9",x"50",x"3A",x"C7",x"E0",x"B7",x"21", -- 0x0FB0
		x"80",x"00",x"28",x"03",x"21",x"80",x"01",x"CD", -- 0x0FB8
		x"67",x"50",x"DD",x"CB",x"0D",x"66",x"28",x"08", -- 0x0FC0
		x"DD",x"7E",x"0F",x"FE",x"E0",x"DA",x"00",x"50", -- 0x0FC8
		x"18",x"04",x"CD",x"E3",x"4F",x"D8",x"CD",x"E8", -- 0x0FD0
		x"2A",x"DD",x"E5",x"E1",x"01",x"2B",x"00",x"09", -- 0x0FD8
		x"C3",x"EF",x"2A",x"DD",x"CB",x"0D",x"66",x"CA", -- 0x0FE0
		x"F5",x"4F",x"DD",x"7E",x"0F",x"FE",x"E0",x"30", -- 0x0FE8
		x"04",x"FE",x"02",x"30",x"0B",x"DD",x"7E",x"0E", -- 0x0FF0
		x"E6",x"FE",x"FE",x"F0",x"28",x"02",x"B7",x"C9", -- 0x0FF8
		x"CD",x"DD",x"66",x"CD",x"CB",x"66",x"37",x"C9", -- 0x1000
		x"21",x"C2",x"B1",x"7E",x"DD",x"77",x"16",x"23", -- 0x1008
		x"7E",x"DD",x"CB",x"02",x"6E",x"28",x"04",x"ED", -- 0x1010
		x"44",x"E6",x"0F",x"DD",x"77",x"19",x"23",x"DD", -- 0x1018
		x"75",x"10",x"DD",x"74",x"11",x"DD",x"7E",x"19", -- 0x1020
		x"07",x"07",x"C6",x"82",x"DD",x"77",x"0C",x"D6", -- 0x1028
		x"02",x"DD",x"77",x"2C",x"C9",x"DD",x"6E",x"10", -- 0x1030
		x"DD",x"66",x"11",x"DD",x"4E",x"24",x"CD",x"BB", -- 0x1038
		x"50",x"DD",x"73",x"24",x"DD",x"7E",x"0F",x"CD", -- 0x1040
		x"AB",x"50",x"DD",x"77",x"0F",x"CD",x"8B",x"50", -- 0x1048
		x"23",x"DD",x"4E",x"25",x"CD",x"BB",x"50",x"DD", -- 0x1050
		x"73",x"25",x"DD",x"7E",x"0E",x"CD",x"A5",x"50", -- 0x1058
		x"DD",x"77",x"0E",x"DD",x"77",x"2E",x"C9",x"DD", -- 0x1060
		x"4E",x"24",x"06",x"00",x"09",x"DD",x"75",x"24", -- 0x1068
		x"DD",x"7E",x"0F",x"84",x"DD",x"77",x"0F",x"57", -- 0x1070
		x"18",x"11",x"DD",x"4E",x"24",x"06",x"00",x"09", -- 0x1078
		x"DD",x"75",x"24",x"DD",x"7E",x"0F",x"94",x"DD", -- 0x1080
		x"77",x"0F",x"57",x"DD",x"7E",x"0D",x"30",x"05", -- 0x1088
		x"EE",x"10",x"DD",x"77",x"0D",x"4F",x"7A",x"C6", -- 0x1090
		x"10",x"DD",x"77",x"2F",x"79",x"30",x"02",x"EE", -- 0x1098
		x"10",x"DD",x"77",x"2D",x"C9",x"DD",x"CB",x"02", -- 0x10A0
		x"6E",x"20",x"06",x"CB",x"46",x"20",x"06",x"18", -- 0x10A8
		x"07",x"CB",x"46",x"20",x"03",x"92",x"18",x"01", -- 0x10B0
		x"82",x"57",x"C9",x"7E",x"E6",x"FC",x"5F",x"16", -- 0x10B8
		x"00",x"42",x"EB",x"29",x"29",x"09",x"EB",x"C9", -- 0x10C0
		x"DD",x"75",x"0F",x"CB",x"44",x"20",x"05",x"DD", -- 0x10C8
		x"CB",x"0D",x"A6",x"C9",x"DD",x"CB",x"0D",x"E6", -- 0x10D0
		x"C9",x"3A",x"46",x"E1",x"4F",x"DD",x"7E",x"0E", -- 0x10D8
		x"C6",x"10",x"57",x"DD",x"7E",x"0F",x"C6",x"08", -- 0x10E0
		x"5F",x"C3",x"F9",x"50",x"DD",x"7E",x"0E",x"C6", -- 0x10E8
		x"08",x"57",x"DD",x"5E",x"0F",x"3A",x"63",x"E1", -- 0x10F0
		x"4F",x"3A",x"C7",x"E0",x"B7",x"C0",x"3A",x"C4", -- 0x10F8
		x"E0",x"B7",x"C0",x"3A",x"C2",x"E0",x"E6",x"02", -- 0x1100
		x"C0",x"21",x"6B",x"E1",x"3A",x"F0",x"E3",x"BE", -- 0x1108
		x"D0",x"DD",x"7E",x"04",x"B7",x"28",x"04",x"DD", -- 0x1110
		x"35",x"04",x"C0",x"DD",x"71",x"04",x"DD",x"7E", -- 0x1118
		x"0D",x"E6",x"10",x"C2",x"F8",x"51",x"DD",x"7E", -- 0x1120
		x"0F",x"4F",x"FE",x"10",x"DA",x"F8",x"51",x"FE", -- 0x1128
		x"EC",x"D2",x"F8",x"51",x"DD",x"7E",x"0E",x"FE", -- 0x1130
		x"10",x"DA",x"F8",x"51",x"FE",x"E0",x"D2",x"F8", -- 0x1138
		x"51",x"3A",x"0E",x"E1",x"C6",x"10",x"6F",x"7A", -- 0x1140
		x"95",x"DC",x"90",x"39",x"FE",x"50",x"D2",x"61", -- 0x1148
		x"51",x"3A",x"0F",x"E1",x"C6",x"08",x"67",x"7B", -- 0x1150
		x"94",x"DC",x"90",x"39",x"FE",x"40",x"DA",x"F8", -- 0x1158
		x"51",x"CD",x"11",x"67",x"DA",x"F8",x"51",x"DD", -- 0x1160
		x"7E",x"01",x"2F",x"E6",x"C0",x"21",x"BE",x"7C", -- 0x1168
		x"20",x"14",x"21",x"DE",x"7C",x"DD",x"CB",x"08", -- 0x1170
		x"7E",x"28",x"0B",x"3A",x"0F",x"E1",x"DD",x"BE", -- 0x1178
		x"0F",x"30",x"03",x"21",x"EE",x"7C",x"DD",x"4E", -- 0x1180
		x"19",x"79",x"FE",x"10",x"38",x"1B",x"FE",x"30", -- 0x1188
		x"38",x"11",x"E6",x"07",x"CA",x"A0",x"51",x"FE", -- 0x1190
		x"04",x"C2",x"F4",x"51",x"79",x"EE",x"14",x"4F", -- 0x1198
		x"79",x"D6",x"20",x"D6",x"10",x"E6",x"18",x"0F", -- 0x11A0
		x"4F",x"CB",x"01",x"06",x"00",x"09",x"DD",x"7E", -- 0x11A8
		x"0F",x"86",x"DD",x"77",x"07",x"23",x"DD",x"7E", -- 0x11B0
		x"0E",x"86",x"DD",x"77",x"06",x"C5",x"CD",x"57", -- 0x11B8
		x"5F",x"51",x"C1",x"DD",x"7E",x"01",x"2F",x"E6", -- 0x11C0
		x"C0",x"20",x"07",x"DD",x"CB",x"08",x"7E",x"C2", -- 0x11C8
		x"E6",x"51",x"21",x"56",x"7C",x"09",x"7E",x"23", -- 0x11D0
		x"66",x"6F",x"7E",x"FE",x"FF",x"28",x"15",x"BB", -- 0x11D8
		x"28",x"04",x"23",x"C3",x"DA",x"51",x"CD",x"86", -- 0x11E0
		x"5E",x"38",x"09",x"21",x"F0",x"E3",x"FD",x"36", -- 0x11E8
		x"00",x"01",x"34",x"C9",x"FD",x"CB",x"00",x"8E", -- 0x11F0
		x"DD",x"36",x"04",x"01",x"37",x"C9",x"CD",x"82", -- 0x11F8
		x"36",x"01",x"01",x"0C",x"16",x"30",x"21",x"09", -- 0x1200
		x"E1",x"CB",x"46",x"20",x"09",x"DD",x"CB",x"02", -- 0x1208
		x"DE",x"01",x"EF",x"04",x"16",x"10",x"DD",x"70", -- 0x1210
		x"19",x"DD",x"71",x"0E",x"DD",x"72",x"0C",x"DD", -- 0x1218
		x"36",x"0F",x"08",x"DD",x"36",x"0D",x"00",x"21", -- 0x1220
		x"A9",x"9F",x"DD",x"75",x"10",x"DD",x"74",x"11", -- 0x1228
		x"7E",x"DD",x"77",x"14",x"DD",x"36",x"18",x"01", -- 0x1230
		x"DD",x"CB",x"00",x"A6",x"DD",x"34",x"03",x"C9", -- 0x1238
		x"CD",x"25",x"34",x"CD",x"25",x"33",x"DD",x"7E", -- 0x1240
		x"18",x"EE",x"01",x"DD",x"77",x"18",x"E6",x"01", -- 0x1248
		x"20",x"08",x"DD",x"7E",x"0D",x"EE",x"01",x"DD", -- 0x1250
		x"77",x"0D",x"CD",x"9A",x"4A",x"D2",x"59",x"3C", -- 0x1258
		x"DD",x"36",x"14",x"FF",x"C3",x"59",x"3C",x"CD", -- 0x1260
		x"E3",x"4A",x"DA",x"87",x"52",x"CD",x"97",x"52", -- 0x1268
		x"DD",x"CB",x"0D",x"66",x"CA",x"E8",x"2A",x"DD", -- 0x1270
		x"7E",x"0F",x"FE",x"F1",x"D2",x"E8",x"2A",x"FE", -- 0x1278
		x"80",x"DA",x"E8",x"2A",x"C3",x"CB",x"66",x"3E", -- 0x1280
		x"BE",x"DD",x"77",x"0C",x"DD",x"36",x"0D",x"0E", -- 0x1288
		x"DD",x"36",x"03",x"04",x"C3",x"70",x"52",x"DD", -- 0x1290
		x"35",x"13",x"C0",x"DD",x"36",x"13",x"02",x"DD", -- 0x1298
		x"7E",x"19",x"DD",x"CB",x"02",x"5E",x"20",x"03", -- 0x12A0
		x"3C",x"18",x"01",x"3D",x"E6",x"0F",x"DD",x"77", -- 0x12A8
		x"19",x"CD",x"0A",x"42",x"DD",x"77",x"0C",x"C9", -- 0x12B0
		x"CD",x"79",x"60",x"D2",x"C5",x"52",x"CD",x"4D", -- 0x12B8
		x"3B",x"D2",x"DE",x"61",x"C9",x"DD",x"CB",x"02", -- 0x12C0
		x"BE",x"21",x"F1",x"52",x"CD",x"D1",x"12",x"CD", -- 0x12C8
		x"55",x"2D",x"DD",x"36",x"0C",x"DE",x"DD",x"36", -- 0x12D0
		x"0D",x"4E",x"DD",x"36",x"16",x"14",x"DD",x"36", -- 0x12D8
		x"03",x"05",x"0E",x"07",x"CD",x"78",x"11",x"C3", -- 0x12E0
		x"E8",x"2A",x"00",x"00",x"00",x"00",x"05",x"00", -- 0x12E8
		x"00",x"00",x"DD",x"35",x"16",x"C0",x"C3",x"CB", -- 0x12F0
		x"66",x"AF",x"32",x"02",x"EC",x"DD",x"77",x"0A", -- 0x12F8
		x"DD",x"77",x"08",x"DD",x"36",x"18",x"00",x"21", -- 0x1300
		x"00",x"00",x"22",x"70",x"E0",x"22",x"72",x"E0", -- 0x1308
		x"22",x"74",x"E0",x"22",x"76",x"E0",x"CD",x"82", -- 0x1310
		x"36",x"CD",x"7B",x"53",x"3A",x"0C",x"E0",x"E6", -- 0x1318
		x"7F",x"C6",x"30",x"6F",x"26",x"00",x"CD",x"AD", -- 0x1320
		x"53",x"21",x"C0",x"01",x"CD",x"C5",x"53",x"21", -- 0x1328
		x"3C",x"06",x"22",x"03",x"EC",x"0E",x"01",x"CD", -- 0x1330
		x"78",x"11",x"CD",x"1A",x"54",x"3A",x"03",x"E1", -- 0x1338
		x"E6",x"3E",x"0F",x"4F",x"06",x"00",x"21",x"FA", -- 0x1340
		x"53",x"09",x"7E",x"32",x"06",x"EC",x"3A",x"0C", -- 0x1348
		x"E0",x"E6",x"03",x"FE",x"03",x"20",x"01",x"AF", -- 0x1350
		x"DD",x"77",x"05",x"21",x"78",x"53",x"4F",x"06", -- 0x1358
		x"00",x"09",x"7E",x"DD",x"77",x"20",x"DD",x"77", -- 0x1360
		x"21",x"DD",x"36",x"04",x"01",x"AF",x"DD",x"77", -- 0x1368
		x"13",x"DD",x"77",x"26",x"DD",x"34",x"03",x"C9", -- 0x1370
		x"01",x"02",x"04",x"21",x"0E",x"7D",x"3A",x"02", -- 0x1378
		x"EC",x"07",x"07",x"07",x"4F",x"06",x"00",x"09", -- 0x1380
		x"7E",x"DD",x"77",x"0C",x"23",x"DD",x"7E",x"0D", -- 0x1388
		x"E6",x"1F",x"B6",x"DD",x"77",x"0D",x"23",x"11", -- 0x1390
		x"12",x"EC",x"CD",x"A0",x"53",x"CD",x"A0",x"53", -- 0x1398
		x"ED",x"A0",x"1A",x"E6",x"1F",x"B6",x"12",x"23", -- 0x13A0
		x"13",x"13",x"13",x"13",x"C9",x"DD",x"77",x"0E", -- 0x13A8
		x"21",x"D2",x"53",x"DD",x"7E",x"0E",x"86",x"32", -- 0x13B0
		x"14",x"EC",x"23",x"86",x"32",x"19",x"EC",x"23", -- 0x13B8
		x"86",x"32",x"1E",x"EC",x"C9",x"DD",x"75",x"0F", -- 0x13C0
		x"CB",x"44",x"20",x"09",x"DD",x"CB",x"0D",x"A6", -- 0x13C8
		x"18",x"07",x"00",x"F0",x"18",x"DD",x"CB",x"0D", -- 0x13D0
		x"E6",x"11",x"13",x"EC",x"01",x"10",x"00",x"CD", -- 0x13D8
		x"E5",x"53",x"CD",x"E5",x"53",x"09",x"1A",x"CB", -- 0x13E0
		x"44",x"20",x"04",x"CB",x"A7",x"18",x"02",x"CB", -- 0x13E8
		x"E7",x"12",x"13",x"13",x"7D",x"12",x"13",x"13", -- 0x13F0
		x"13",x"C9",x"88",x"80",x"70",x"88",x"88",x"78", -- 0x13F8
		x"68",x"88",x"88",x"58",x"70",x"88",x"78",x"68", -- 0x1400
		x"58",x"88",x"78",x"60",x"50",x"88",x"70",x"60", -- 0x1408
		x"50",x"88",x"68",x"60",x"50",x"88",x"50",x"40", -- 0x1410
		x"30",x"88",x"CD",x"E8",x"2A",x"21",x"11",x"EC", -- 0x1418
		x"CD",x"26",x"54",x"CD",x"26",x"54",x"5E",x"16", -- 0x1420
		x"EB",x"23",x"01",x"04",x"00",x"ED",x"B0",x"C9", -- 0x1428
		x"01",x"01",x"00",x"CD",x"09",x"62",x"09",x"CD", -- 0x1430
		x"C5",x"53",x"CD",x"1A",x"54",x"3A",x"1D",x"EC", -- 0x1438
		x"DD",x"B6",x"0D",x"E6",x"10",x"C0",x"DD",x"34", -- 0x1440
		x"03",x"AF",x"DD",x"77",x"14",x"DD",x"77",x"15", -- 0x1448
		x"C9",x"DD",x"7E",x"13",x"CD",x"F7",x"66",x"67", -- 0x1450
		x"54",x"AD",x"54",x"F3",x"54",x"78",x"55",x"A6", -- 0x1458
		x"55",x"CD",x"55",x"35",x"56",x"9D",x"56",x"CD", -- 0x1460
		x"9C",x"55",x"CD",x"CA",x"56",x"3A",x"06",x"EC", -- 0x1468
		x"DD",x"BE",x"0F",x"D2",x"1A",x"54",x"DD",x"7E", -- 0x1470
		x"0E",x"FE",x"70",x"3E",x"09",x"38",x"01",x"3C", -- 0x1478
		x"DD",x"77",x"15",x"DD",x"CB",x"01",x"FE",x"21", -- 0x1480
		x"CE",x"7D",x"11",x"DB",x"7D",x"7E",x"DD",x"77", -- 0x1488
		x"14",x"23",x"DD",x"75",x"10",x"DD",x"74",x"11", -- 0x1490
		x"1A",x"DD",x"77",x"17",x"13",x"DD",x"73",x"1E", -- 0x1498
		x"DD",x"72",x"1F",x"DD",x"34",x"13",x"DD",x"CB", -- 0x14A0
		x"00",x"A6",x"C3",x"1A",x"54",x"CD",x"9C",x"55", -- 0x14A8
		x"CD",x"F2",x"56",x"DD",x"7E",x"0E",x"DD",x"CB", -- 0x14B0
		x"15",x"46",x"20",x"06",x"FE",x"48",x"30",x"17", -- 0x14B8
		x"18",x"04",x"FE",x"98",x"38",x"11",x"21",x"E8", -- 0x14C0
		x"7D",x"11",x"F3",x"7D",x"DD",x"7E",x"15",x"EE", -- 0x14C8
		x"0C",x"DD",x"77",x"15",x"C3",x"8D",x"54",x"CD", -- 0x14D0
		x"D5",x"58",x"DD",x"35",x"14",x"C2",x"E5",x"54", -- 0x14D8
		x"0E",x"01",x"CD",x"46",x"55",x"DD",x"35",x"17", -- 0x14E0
		x"C2",x"1A",x"54",x"0E",x"01",x"CD",x"5E",x"55", -- 0x14E8
		x"C3",x"1A",x"54",x"CD",x"9C",x"55",x"CD",x"F2", -- 0x14F0
		x"56",x"CD",x"D5",x"58",x"DD",x"35",x"14",x"20", -- 0x14F8
		x"05",x"0E",x"01",x"CD",x"46",x"55",x"3A",x"C7", -- 0x1500
		x"E0",x"B7",x"28",x"07",x"DD",x"36",x"13",x"04", -- 0x1508
		x"C3",x"1A",x"54",x"DD",x"35",x"17",x"C2",x"1A", -- 0x1510
		x"54",x"CD",x"5E",x"55",x"C2",x"1A",x"54",x"DD", -- 0x1518
		x"7E",x"15",x"EE",x"03",x"DD",x"77",x"15",x"CD", -- 0x1520
		x"2D",x"55",x"C3",x"8D",x"54",x"21",x"0C",x"7E", -- 0x1528
		x"DD",x"7E",x"05",x"07",x"CD",x"3D",x"55",x"23", -- 0x1530
		x"7E",x"23",x"66",x"6F",x"C9",x"07",x"4F",x"06", -- 0x1538
		x"00",x"09",x"5E",x"23",x"56",x"C9",x"DD",x"6E", -- 0x1540
		x"10",x"DD",x"66",x"11",x"23",x"7E",x"B7",x"DD", -- 0x1548
		x"71",x"14",x"C8",x"DD",x"77",x"14",x"23",x"DD", -- 0x1550
		x"75",x"10",x"DD",x"74",x"11",x"C9",x"DD",x"6E", -- 0x1558
		x"1E",x"DD",x"66",x"1F",x"23",x"7E",x"B7",x"DD", -- 0x1560
		x"71",x"17",x"CA",x"1A",x"54",x"DD",x"77",x"17", -- 0x1568
		x"23",x"DD",x"75",x"1E",x"DD",x"74",x"1F",x"C9", -- 0x1570
		x"CD",x"9C",x"55",x"CD",x"F2",x"56",x"CD",x"7C", -- 0x1578
		x"58",x"3A",x"C7",x"E0",x"B7",x"20",x"0B",x"2A", -- 0x1580
		x"03",x"EC",x"2D",x"20",x"09",x"2E",x"3C",x"25", -- 0x1588
		x"20",x"04",x"DD",x"36",x"13",x"04",x"22",x"03", -- 0x1590
		x"EC",x"C3",x"1A",x"54",x"3A",x"C7",x"E0",x"B7", -- 0x1598
		x"C8",x"DD",x"36",x"13",x"04",x"C9",x"CD",x"09", -- 0x15A0
		x"62",x"01",x"01",x"00",x"09",x"CD",x"C5",x"53", -- 0x15A8
		x"CD",x"1A",x"54",x"DD",x"CB",x"0D",x"66",x"C8", -- 0x15B0
		x"DD",x"7E",x"0F",x"FE",x"C0",x"D0",x"CD",x"B3", -- 0x15B8
		x"56",x"AF",x"DD",x"77",x"00",x"32",x"05",x"EC", -- 0x15C0
		x"0E",x"0B",x"C3",x"78",x"11",x"DD",x"35",x"16", -- 0x15C8
		x"20",x"16",x"21",x"02",x"EC",x"34",x"7E",x"FE", -- 0x15D0
		x"07",x"30",x"16",x"DD",x"36",x"16",x"08",x"CD", -- 0x15D8
		x"7B",x"53",x"DD",x"7E",x"0E",x"CD",x"AD",x"53", -- 0x15E0
		x"21",x"00",x"01",x"CD",x"01",x"59",x"C3",x"B0", -- 0x15E8
		x"55",x"DD",x"34",x"13",x"DD",x"36",x"16",x"07", -- 0x15F0
		x"AF",x"DD",x"77",x"1C",x"6F",x"67",x"22",x"1D", -- 0x15F8
		x"EC",x"CD",x"29",x"56",x"DD",x"7E",x"1A",x"C6", -- 0x1600
		x"06",x"4F",x"3A",x"13",x"EC",x"E6",x"10",x"F6", -- 0x1608
		x"60",x"B1",x"32",x"13",x"EC",x"3A",x"18",x"EC", -- 0x1610
		x"E6",x"10",x"F6",x"60",x"B1",x"32",x"18",x"EC", -- 0x1618
		x"3A",x"14",x"EC",x"32",x"19",x"EC",x"C3",x"1A", -- 0x1620
		x"54",x"CD",x"2E",x"64",x"32",x"17",x"EC",x"23", -- 0x1628
		x"7E",x"32",x"12",x"EC",x"C9",x"DD",x"35",x"16", -- 0x1630
		x"C2",x"1A",x"54",x"DD",x"7E",x"1C",x"3C",x"FE", -- 0x1638
		x"0A",x"30",x"0D",x"DD",x"77",x"1C",x"CD",x"29", -- 0x1640
		x"56",x"DD",x"36",x"16",x"07",x"C3",x"1A",x"54", -- 0x1648
		x"3A",x"07",x"EC",x"07",x"07",x"4F",x"06",x"00", -- 0x1650
		x"21",x"8C",x"7E",x"09",x"7E",x"32",x"12",x"EC", -- 0x1658
		x"23",x"7E",x"DD",x"77",x"0C",x"3A",x"13",x"EC", -- 0x1660
		x"E6",x"10",x"F6",x"0E",x"32",x"13",x"EC",x"DD", -- 0x1668
		x"77",x"0D",x"3A",x"14",x"EC",x"C6",x"10",x"DD", -- 0x1670
		x"77",x"0E",x"3A",x"15",x"EC",x"DD",x"77",x"0F", -- 0x1678
		x"DD",x"36",x"16",x"40",x"21",x"00",x"00",x"22", -- 0x1680
		x"18",x"EC",x"3A",x"07",x"EC",x"3C",x"FE",x"0E", -- 0x1688
		x"38",x"02",x"3E",x"0E",x"32",x"07",x"EC",x"DD", -- 0x1690
		x"34",x"13",x"C3",x"1A",x"54",x"DD",x"35",x"16", -- 0x1698
		x"C0",x"AF",x"6F",x"67",x"DD",x"77",x"0D",x"DD", -- 0x16A0
		x"77",x"0E",x"22",x"13",x"EC",x"CD",x"1A",x"54", -- 0x16A8
		x"C3",x"BE",x"55",x"CD",x"02",x"67",x"11",x"11", -- 0x16B0
		x"EC",x"01",x"05",x"00",x"CD",x"C2",x"56",x"CD", -- 0x16B8
		x"C2",x"56",x"1A",x"CD",x"05",x"67",x"EB",x"09", -- 0x16C0
		x"EB",x"C9",x"01",x"01",x"00",x"CD",x"09",x"62", -- 0x16C8
		x"09",x"C3",x"C5",x"53",x"3A",x"00",x"E0",x"07", -- 0x16D0
		x"D2",x"EC",x"56",x"DD",x"E5",x"E1",x"29",x"29", -- 0x16D8
		x"29",x"7C",x"E6",x"0F",x"21",x"E0",x"E0",x"85", -- 0x16E0
		x"6F",x"34",x"7E",x"C9",x"21",x"2D",x"E0",x"34", -- 0x16E8
		x"7E",x"C9",x"3A",x"C4",x"E0",x"B7",x"C0",x"3A", -- 0x16F0
		x"C7",x"E0",x"B7",x"C0",x"3A",x"C2",x"E0",x"E6", -- 0x16F8
		x"02",x"C0",x"3A",x"44",x"E1",x"B7",x"C0",x"DD", -- 0x1700
		x"CB",x"26",x"4E",x"CA",x"18",x"57",x"DD",x"35", -- 0x1708
		x"27",x"C0",x"DD",x"7E",x"28",x"C3",x"83",x"57", -- 0x1710
		x"DD",x"35",x"04",x"C0",x"DD",x"36",x"04",x"01", -- 0x1718
		x"2A",x"0E",x"E1",x"DD",x"56",x"0E",x"DD",x"5E", -- 0x1720
		x"0F",x"7B",x"C6",x"18",x"94",x"DC",x"90",x"39", -- 0x1728
		x"FE",x"48",x"30",x"08",x"7A",x"95",x"DC",x"90", -- 0x1730
		x"39",x"FE",x"40",x"D8",x"7B",x"BC",x"30",x"12", -- 0x1738
		x"C6",x"30",x"5F",x"BC",x"DA",x"52",x"57",x"7A", -- 0x1740
		x"BD",x"3E",x"01",x"D2",x"7D",x"57",x"3C",x"C3", -- 0x1748
		x"7D",x"57",x"0E",x"00",x"7D",x"92",x"30",x"04", -- 0x1750
		x"ED",x"44",x"0E",x"04",x"47",x"7C",x"93",x"30", -- 0x1758
		x"04",x"ED",x"44",x"CB",x"C9",x"B8",x"30",x"01", -- 0x1760
		x"0C",x"06",x"00",x"21",x"47",x"58",x"09",x"3A", -- 0x1768
		x"EF",x"E0",x"3C",x"32",x"EF",x"E0",x"E6",x"04", -- 0x1770
		x"7E",x"28",x"02",x"0F",x"0F",x"E6",x"03",x"07", -- 0x1778
		x"DD",x"77",x"28",x"4F",x"06",x"00",x"21",x"76", -- 0x1780
		x"7D",x"09",x"7E",x"DD",x"86",x"0F",x"DA",x"FC", -- 0x1788
		x"57",x"DD",x"77",x"07",x"23",x"7E",x"DD",x"86", -- 0x1790
		x"0E",x"38",x"61",x"DD",x"77",x"06",x"CD",x"11", -- 0x1798
		x"67",x"DA",x"FC",x"57",x"DD",x"CB",x"26",x"4E", -- 0x17A0
		x"C2",x"E9",x"57",x"CD",x"D4",x"5D",x"DA",x"F8", -- 0x17A8
		x"57",x"FD",x"E5",x"E1",x"CD",x"EB",x"2A",x"FD", -- 0x17B0
		x"36",x"00",x"01",x"CD",x"0F",x"58",x"DD",x"7E", -- 0x17B8
		x"29",x"86",x"DD",x"CB",x"26",x"46",x"28",x"02", -- 0x17C0
		x"96",x"96",x"DD",x"77",x"29",x"21",x"F0",x"E3", -- 0x17C8
		x"34",x"DD",x"7E",x"26",x"C6",x"20",x"30",x"01", -- 0x17D0
		x"AF",x"DD",x"77",x"26",x"3A",x"78",x"E1",x"DD", -- 0x17D8
		x"77",x"04",x"3A",x"79",x"E1",x"DD",x"77",x"27", -- 0x17E0
		x"C9",x"DD",x"7E",x"29",x"CD",x"05",x"58",x"5E", -- 0x17E8
		x"DD",x"56",x"2A",x"CD",x"86",x"5E",x"18",x"B6", -- 0x17F0
		x"FD",x"36",x"00",x"00",x"DD",x"36",x"04",x"01", -- 0x17F8
		x"DD",x"36",x"27",x"01",x"C9",x"21",x"47",x"5F", -- 0x1800
		x"E6",x"0F",x"4F",x"06",x"00",x"09",x"C9",x"3A", -- 0x1808
		x"03",x"E1",x"4F",x"E6",x"03",x"FE",x"03",x"28", -- 0x1810
		x"21",x"3A",x"04",x"C0",x"07",x"07",x"07",x"07", -- 0x1818
		x"E6",x"06",x"4F",x"06",x"00",x"21",x"4F",x"58", -- 0x1820
		x"09",x"7E",x"23",x"66",x"6F",x"3A",x"03",x"E1", -- 0x1828
		x"BE",x"38",x"01",x"7E",x"23",x"4F",x"06",x"00", -- 0x1830
		x"09",x"C9",x"79",x"0F",x"0F",x"E6",x"07",x"4F", -- 0x1838
		x"06",x"00",x"21",x"74",x"58",x"09",x"C9",x"00", -- 0x1840
		x"02",x"0B",x"0A",x"00",x"01",x"07",x"05",x"72", -- 0x1848
		x"58",x"72",x"58",x"57",x"58",x"6A",x"58",x"11", -- 0x1850
		x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x1858
		x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02", -- 0x1860
		x"02",x"01",x"06",x"02",x"02",x"02",x"01",x"02", -- 0x1868
		x"02",x"01",x"00",x"01",x"02",x"02",x"01",x"02", -- 0x1870
		x"02",x"01",x"01",x"02",x"CD",x"D5",x"58",x"DD", -- 0x1878
		x"35",x"14",x"20",x"2C",x"CD",x"46",x"55",x"20", -- 0x1880
		x"27",x"21",x"00",x"7E",x"DD",x"7E",x"05",x"CD", -- 0x1888
		x"3D",x"55",x"1A",x"DD",x"77",x"14",x"13",x"DD", -- 0x1890
		x"73",x"10",x"DD",x"72",x"11",x"DD",x"35",x"21", -- 0x1898
		x"20",x"0E",x"DD",x"7E",x"20",x"DD",x"77",x"21", -- 0x18A0
		x"DD",x"7E",x"15",x"EE",x"03",x"DD",x"77",x"15", -- 0x18A8
		x"DD",x"35",x"17",x"C0",x"CD",x"5E",x"55",x"C0", -- 0x18B0
		x"21",x"06",x"7E",x"DD",x"7E",x"05",x"CD",x"3D", -- 0x18B8
		x"55",x"1A",x"DD",x"77",x"17",x"13",x"DD",x"73", -- 0x18C0
		x"1E",x"DD",x"72",x"1F",x"DD",x"7E",x"15",x"EE", -- 0x18C8
		x"0C",x"DD",x"77",x"15",x"C9",x"DD",x"6E",x"10", -- 0x18D0
		x"DD",x"66",x"11",x"6E",x"26",x"00",x"44",x"29", -- 0x18D8
		x"DD",x"4E",x"25",x"09",x"DD",x"75",x"25",x"DD", -- 0x18E0
		x"CB",x"15",x"4E",x"DD",x"7E",x"0E",x"20",x"03", -- 0x18E8
		x"84",x"18",x"01",x"94",x"CD",x"AD",x"53",x"DD", -- 0x18F0
		x"6E",x"1E",x"DD",x"66",x"1F",x"6E",x"26",x"00", -- 0x18F8
		x"29",x"DD",x"4E",x"24",x"06",x"00",x"09",x"DD", -- 0x1900
		x"75",x"24",x"DD",x"CB",x"15",x"56",x"DD",x"7E", -- 0x1908
		x"0F",x"20",x"03",x"84",x"18",x"01",x"94",x"DD", -- 0x1910
		x"77",x"0F",x"6F",x"26",x"00",x"30",x"08",x"DD", -- 0x1918
		x"CB",x"0D",x"66",x"20",x"09",x"18",x"06",x"DD", -- 0x1920
		x"CB",x"0D",x"66",x"28",x"01",x"24",x"C3",x"C5", -- 0x1928
		x"53",x"3E",x"01",x"32",x"B4",x"E7",x"21",x"E8", -- 0x1930
		x"7E",x"0E",x"10",x"3A",x"03",x"E1",x"FE",x"1E", -- 0x1938
		x"38",x"02",x"0E",x"12",x"11",x"40",x"EB",x"06", -- 0x1940
		x"10",x"C5",x"ED",x"A0",x"C1",x"7E",x"E6",x"E0", -- 0x1948
		x"B1",x"12",x"23",x"13",x"13",x"13",x"10",x"F1", -- 0x1950
		x"21",x"71",x"80",x"DD",x"CB",x"01",x"4E",x"20", -- 0x1958
		x"02",x"26",x"00",x"DD",x"75",x"0E",x"DD",x"74", -- 0x1960
		x"0F",x"DD",x"75",x"1E",x"DD",x"74",x"1F",x"DD", -- 0x1968
		x"7E",x"1A",x"F6",x"30",x"DD",x"77",x"20",x"DD", -- 0x1970
		x"77",x"0D",x"CD",x"4F",x"5D",x"AF",x"DD",x"77", -- 0x1978
		x"24",x"DD",x"CB",x"01",x"4E",x"21",x"08",x"7F", -- 0x1980
		x"20",x"03",x"21",x"11",x"7F",x"CD",x"2B",x"5D", -- 0x1988
		x"3E",x"01",x"DD",x"77",x"04",x"32",x"DE",x"E9", -- 0x1990
		x"3C",x"32",x"E6",x"E9",x"3A",x"0C",x"E0",x"E6", -- 0x1998
		x"07",x"3C",x"32",x"D4",x"E9",x"21",x"E0",x"E0", -- 0x19A0
		x"86",x"77",x"E6",x"07",x"3C",x"32",x"DC",x"E9", -- 0x19A8
		x"23",x"86",x"77",x"E6",x"07",x"3C",x"32",x"E4", -- 0x19B0
		x"E9",x"AF",x"67",x"6F",x"32",x"D6",x"E9",x"DD", -- 0x19B8
		x"77",x"1C",x"DD",x"77",x"26",x"32",x"D0",x"E9", -- 0x19C0
		x"32",x"D8",x"E9",x"32",x"E0",x"E9",x"32",x"F8", -- 0x19C8
		x"E9",x"22",x"F9",x"E9",x"DD",x"77",x"13",x"0E", -- 0x19D0
		x"01",x"CD",x"78",x"11",x"0E",x"10",x"CD",x"78", -- 0x19D8
		x"11",x"0E",x"1A",x"CD",x"78",x"11",x"21",x"E0", -- 0x19E0
		x"00",x"DD",x"75",x"22",x"DD",x"74",x"23",x"DD", -- 0x19E8
		x"36",x"03",x"01",x"C9",x"DD",x"6E",x"22",x"DD", -- 0x19F0
		x"66",x"23",x"7D",x"B4",x"28",x"10",x"2B",x"DD", -- 0x19F8
		x"75",x"22",x"DD",x"74",x"23",x"7D",x"B4",x"20", -- 0x1A00
		x"05",x"0E",x"14",x"CD",x"78",x"11",x"DD",x"7E", -- 0x1A08
		x"13",x"E6",x"01",x"CD",x"F7",x"66",x"1A",x"5A", -- 0x1A10
		x"30",x"5A",x"CD",x"A6",x"5C",x"CD",x"FB",x"5C", -- 0x1A18
		x"3A",x"41",x"EB",x"CB",x"67",x"C0",x"3A",x"43", -- 0x1A20
		x"EB",x"FE",x"40",x"D8",x"DD",x"34",x"13",x"C9", -- 0x1A28
		x"CD",x"A6",x"5C",x"CD",x"D0",x"5B",x"CD",x"D3", -- 0x1A30
		x"5A",x"C3",x"FB",x"5C",x"DD",x"7E",x"13",x"CD", -- 0x1A38
		x"F7",x"66",x"46",x"5A",x"6E",x"5A",x"DD",x"35", -- 0x1A40
		x"14",x"C0",x"AF",x"67",x"6F",x"22",x"51",x"EB", -- 0x1A48
		x"22",x"55",x"EB",x"22",x"59",x"EB",x"22",x"71", -- 0x1A50
		x"EB",x"22",x"75",x"EB",x"22",x"79",x"EB",x"3A", -- 0x1A58
		x"03",x"E1",x"E6",x"18",x"FE",x"18",x"C2",x"BC", -- 0x1A60
		x"5A",x"DD",x"36",x"13",x"01",x"C9",x"DD",x"E5", -- 0x1A68
		x"DD",x"21",x"05",x"A2",x"CD",x"CC",x"2C",x"DD", -- 0x1A70
		x"E1",x"21",x"F2",x"D0",x"CD",x"C1",x"5A",x"21", -- 0x1A78
		x"F6",x"D0",x"CD",x"C1",x"5A",x"21",x"F2",x"D0", -- 0x1A80
		x"CD",x"C7",x"5A",x"21",x"12",x"D3",x"CD",x"C7", -- 0x1A88
		x"5A",x"21",x"34",x"D1",x"11",x"76",x"A6",x"06", -- 0x1A90
		x"0E",x"CD",x"EE",x"01",x"06",x"1E",x"DF",x"21", -- 0x1A98
		x"DC",x"A6",x"CD",x"22",x"02",x"06",x"1E",x"DF", -- 0x1AA0
		x"21",x"FE",x"A6",x"CD",x"22",x"02",x"06",x"82", -- 0x1AA8
		x"DF",x"21",x"41",x"D0",x"01",x"1D",x"1C",x"16", -- 0x1AB0
		x"30",x"CD",x"53",x"02",x"DD",x"36",x"00",x"00", -- 0x1AB8
		x"C9",x"01",x"31",x"12",x"C3",x"49",x"02",x"01", -- 0x1AC0
		x"04",x"00",x"16",x"31",x"C3",x"E2",x"01",x"D0", -- 0x1AC8
		x"86",x"4C",x"44",x"3A",x"C4",x"E0",x"B7",x"C0", -- 0x1AD0
		x"DD",x"CB",x"26",x"4E",x"CA",x"E9",x"5A",x"DD", -- 0x1AD8
		x"35",x"27",x"C0",x"DD",x"7E",x"28",x"C3",x"45", -- 0x1AE0
		x"5B",x"DD",x"35",x"04",x"C0",x"DD",x"36",x"04", -- 0x1AE8
		x"01",x"2A",x"0E",x"E1",x"DD",x"56",x"0E",x"DD", -- 0x1AF0
		x"7E",x"0F",x"C6",x"08",x"5F",x"BC",x"30",x"14", -- 0x1AF8
		x"C6",x"5C",x"5F",x"BC",x"DA",x"14",x"5B",x"7A", -- 0x1B00
		x"C6",x"10",x"BD",x"3E",x"01",x"D2",x"3F",x"5B", -- 0x1B08
		x"3C",x"C3",x"3F",x"5B",x"0E",x"00",x"7D",x"92", -- 0x1B10
		x"30",x"04",x"ED",x"44",x"0E",x"04",x"47",x"7C", -- 0x1B18
		x"93",x"30",x"04",x"ED",x"44",x"CB",x"C9",x"B8", -- 0x1B20
		x"30",x"01",x"0C",x"06",x"00",x"21",x"C8",x"5B", -- 0x1B28
		x"09",x"3A",x"EF",x"E0",x"3C",x"32",x"EF",x"E0", -- 0x1B30
		x"E6",x"04",x"7E",x"28",x"02",x"0F",x"0F",x"E6", -- 0x1B38
		x"03",x"07",x"DD",x"77",x"28",x"4F",x"06",x"00", -- 0x1B40
		x"21",x"28",x"7F",x"09",x"7E",x"DD",x"86",x"0F", -- 0x1B48
		x"DA",x"BF",x"5B",x"DD",x"77",x"07",x"23",x"7E", -- 0x1B50
		x"DD",x"86",x"0E",x"DD",x"77",x"06",x"CD",x"11", -- 0x1B58
		x"67",x"DA",x"BF",x"5B",x"DD",x"CB",x"26",x"4E", -- 0x1B60
		x"C2",x"AC",x"5B",x"CD",x"57",x"5F",x"51",x"3E", -- 0x1B68
		x"A2",x"CD",x"E3",x"5D",x"DA",x"BB",x"5B",x"FD", -- 0x1B70
		x"E5",x"E1",x"CD",x"EB",x"2A",x"FD",x"36",x"00", -- 0x1B78
		x"01",x"DD",x"7E",x"29",x"3C",x"DD",x"CB",x"26", -- 0x1B80
		x"46",x"28",x"02",x"D6",x"02",x"DD",x"77",x"29", -- 0x1B88
		x"21",x"F0",x"E3",x"34",x"DD",x"7E",x"26",x"C6", -- 0x1B90
		x"20",x"30",x"01",x"AF",x"DD",x"77",x"26",x"3A", -- 0x1B98
		x"F0",x"E9",x"DD",x"77",x"04",x"3A",x"F1",x"E9", -- 0x1BA0
		x"DD",x"77",x"27",x"C9",x"DD",x"7E",x"29",x"CD", -- 0x1BA8
		x"05",x"58",x"5E",x"DD",x"56",x"2A",x"CD",x"86", -- 0x1BB0
		x"5E",x"18",x"B9",x"FD",x"36",x"00",x"00",x"DD", -- 0x1BB8
		x"36",x"04",x"01",x"DD",x"36",x"27",x"01",x"C9", -- 0x1BC0
		x"00",x"02",x"0B",x"0A",x"00",x"01",x"07",x"05", -- 0x1BC8
		x"21",x"D0",x"E9",x"22",x"FC",x"E9",x"CD",x"E8", -- 0x1BD0
		x"5B",x"21",x"D8",x"E9",x"22",x"FC",x"E9",x"CD", -- 0x1BD8
		x"E8",x"5B",x"21",x"E0",x"E9",x"22",x"FC",x"E9", -- 0x1BE0
		x"3A",x"C4",x"E0",x"B7",x"C0",x"2A",x"FC",x"E9", -- 0x1BE8
		x"E5",x"FD",x"E1",x"CB",x"4E",x"CA",x"FF",x"5B", -- 0x1BF0
		x"FD",x"35",x"01",x"C0",x"C3",x"07",x"5C",x"FD", -- 0x1BF8
		x"35",x"04",x"C0",x"FD",x"36",x"04",x"01",x"21", -- 0x1C00
		x"32",x"7F",x"FD",x"7E",x"06",x"B7",x"28",x"09", -- 0x1C08
		x"21",x"30",x"7F",x"3D",x"28",x"03",x"21",x"34", -- 0x1C10
		x"7F",x"7E",x"DD",x"86",x"0F",x"DA",x"97",x"5C", -- 0x1C18
		x"DD",x"77",x"07",x"23",x"7E",x"DD",x"86",x"0E", -- 0x1C20
		x"DD",x"77",x"06",x"CD",x"11",x"67",x"DA",x"97", -- 0x1C28
		x"5C",x"2A",x"FC",x"E9",x"CB",x"4E",x"C2",x"79", -- 0x1C30
		x"5C",x"CD",x"8E",x"5D",x"DA",x"93",x"5C",x"FD", -- 0x1C38
		x"E5",x"E1",x"CD",x"EB",x"2A",x"FD",x"36",x"00", -- 0x1C40
		x"01",x"2A",x"FC",x"E9",x"E5",x"FD",x"E1",x"46", -- 0x1C48
		x"FD",x"7E",x"02",x"3C",x"CB",x"40",x"28",x"02", -- 0x1C50
		x"D6",x"02",x"FD",x"77",x"02",x"21",x"F0",x"E3", -- 0x1C58
		x"34",x"FD",x"7E",x"00",x"C6",x"20",x"30",x"01", -- 0x1C60
		x"AF",x"FD",x"77",x"00",x"3A",x"F0",x"E9",x"FD", -- 0x1C68
		x"77",x"04",x"3A",x"F1",x"E9",x"FD",x"77",x"01", -- 0x1C70
		x"C9",x"FD",x"E5",x"2A",x"FC",x"E9",x"E5",x"FD", -- 0x1C78
		x"E1",x"FD",x"7E",x"02",x"CD",x"05",x"58",x"5E", -- 0x1C80
		x"FD",x"7E",x"03",x"57",x"FD",x"E1",x"CD",x"86", -- 0x1C88
		x"5E",x"18",x"A9",x"FD",x"36",x"00",x"00",x"2A", -- 0x1C90
		x"FC",x"E9",x"E5",x"FD",x"E1",x"3E",x"01",x"FD", -- 0x1C98
		x"77",x"04",x"FD",x"77",x"01",x"C9",x"3A",x"F8", -- 0x1CA0
		x"E9",x"B7",x"C8",x"07",x"4F",x"06",x"00",x"21", -- 0x1CA8
		x"F5",x"5C",x"09",x"3A",x"F9",x"E9",x"B7",x"28", -- 0x1CB0
		x"05",x"3D",x"32",x"F9",x"E9",x"C0",x"3A",x"FA", -- 0x1CB8
		x"E9",x"EE",x"01",x"32",x"FA",x"E9",x"E6",x"01", -- 0x1CC0
		x"4F",x"20",x"01",x"23",x"7E",x"32",x"F9",x"E9", -- 0x1CC8
		x"CB",x"41",x"DD",x"7E",x"1A",x"20",x"02",x"EE", -- 0x1CD0
		x"02",x"4F",x"DD",x"7E",x"20",x"E6",x"F0",x"B1", -- 0x1CD8
		x"DD",x"77",x"20",x"DD",x"77",x"0D",x"21",x"41", -- 0x1CE0
		x"EB",x"11",x"04",x"00",x"06",x"10",x"7E",x"E6", -- 0x1CE8
		x"F0",x"B1",x"77",x"19",x"10",x"F8",x"C9",x"08", -- 0x1CF0
		x"04",x"04",x"03",x"DD",x"6E",x"10",x"DD",x"66", -- 0x1CF8
		x"11",x"E5",x"DD",x"4E",x"24",x"CD",x"BB",x"50", -- 0x1D00
		x"DD",x"73",x"24",x"DD",x"7E",x"0F",x"CD",x"AB", -- 0x1D08
		x"50",x"DD",x"77",x"0F",x"DD",x"77",x"1F",x"DD", -- 0x1D10
		x"7E",x"0D",x"30",x"05",x"EE",x"10",x"DD",x"77", -- 0x1D18
		x"0D",x"DD",x"77",x"20",x"E1",x"DD",x"35",x"12", -- 0x1D20
		x"20",x"25",x"23",x"7E",x"B7",x"28",x"0C",x"DD", -- 0x1D28
		x"77",x"12",x"23",x"DD",x"75",x"10",x"DD",x"74", -- 0x1D30
		x"11",x"18",x"14",x"DD",x"7E",x"01",x"EE",x"02", -- 0x1D38
		x"DD",x"77",x"01",x"21",x"16",x"7F",x"E6",x"02", -- 0x1D40
		x"28",x"E1",x"21",x"1F",x"7F",x"18",x"DC",x"DD", -- 0x1D48
		x"7E",x"20",x"4F",x"21",x"C8",x"7E",x"06",x"10", -- 0x1D50
		x"FD",x"21",x"40",x"EB",x"DD",x"7E",x"1E",x"86", -- 0x1D58
		x"FD",x"77",x"02",x"23",x"DD",x"7E",x"1F",x"86", -- 0x1D60
		x"FD",x"77",x"03",x"30",x"0F",x"79",x"EE",x"10", -- 0x1D68
		x"5F",x"FD",x"7E",x"01",x"E6",x"E3",x"B3",x"FD", -- 0x1D70
		x"77",x"01",x"18",x"09",x"FD",x"7E",x"01",x"E6", -- 0x1D78
		x"E3",x"B1",x"FD",x"77",x"01",x"23",x"11",x"04", -- 0x1D80
		x"00",x"FD",x"19",x"10",x"CF",x"C9",x"FD",x"E5", -- 0x1D88
		x"CD",x"57",x"5F",x"2A",x"FC",x"E9",x"E5",x"FD", -- 0x1D90
		x"E1",x"3E",x"A2",x"FD",x"77",x"00",x"51",x"06", -- 0x1D98
		x"00",x"21",x"47",x"5F",x"7B",x"BE",x"28",x"04", -- 0x1DA0
		x"04",x"23",x"18",x"F9",x"78",x"FD",x"77",x"02", -- 0x1DA8
		x"3A",x"F0",x"E0",x"0F",x"38",x"0D",x"FD",x"7E", -- 0x1DB0
		x"00",x"F6",x"01",x"FD",x"77",x"00",x"78",x"C6", -- 0x1DB8
		x"01",x"18",x"03",x"78",x"D6",x"01",x"E6",x"0F", -- 0x1DC0
		x"FD",x"77",x"02",x"CD",x"05",x"58",x"5E",x"FD", -- 0x1DC8
		x"E1",x"C3",x"86",x"5E",x"CD",x"57",x"5F",x"51", -- 0x1DD0
		x"CD",x"0F",x"58",x"7E",x"3D",x"3E",x"A2",x"20", -- 0x1DD8
		x"02",x"3E",x"62",x"DD",x"77",x"26",x"06",x"00", -- 0x1DE0
		x"21",x"47",x"5F",x"7B",x"BE",x"28",x"04",x"04", -- 0x1DE8
		x"23",x"18",x"F9",x"DD",x"70",x"29",x"DD",x"7E", -- 0x1DF0
		x"28",x"B7",x"EA",x"2B",x"5E",x"FE",x"02",x"78", -- 0x1DF8
		x"28",x"15",x"DD",x"CB",x"26",x"C6",x"FE",x"07", -- 0x1E00
		x"38",x"04",x"3E",x"07",x"18",x"06",x"FE",x"03", -- 0x1E08
		x"30",x"02",x"3E",x"03",x"3C",x"18",x"66",x"B7", -- 0x1E10
		x"28",x"0E",x"FE",x"09",x"30",x"04",x"3E",x"09", -- 0x1E18
		x"18",x"06",x"FE",x"0D",x"30",x"02",x"3E",x"0D", -- 0x1E20
		x"3D",x"18",x"52",x"28",x"25",x"3A",x"0C",x"E0", -- 0x1E28
		x"07",x"78",x"30",x"0C",x"FE",x"0E",x"30",x"2F", -- 0x1E30
		x"FE",x"04",x"38",x"2B",x"3E",x"04",x"18",x"27", -- 0x1E38
		x"FE",x"0C",x"30",x"38",x"FE",x"02",x"38",x"34", -- 0x1E40
		x"FE",x"08",x"3E",x"02",x"38",x"2E",x"3E",x"0C", -- 0x1E48
		x"18",x"2A",x"3A",x"0C",x"E0",x"07",x"78",x"30", -- 0x1E50
		x"15",x"FE",x"06",x"30",x"04",x"3E",x"06",x"18", -- 0x1E58
		x"06",x"FE",x"0C",x"38",x"02",x"3E",x"0C",x"DD", -- 0x1E60
		x"CB",x"26",x"C6",x"3C",x"18",x"0F",x"FE",x"04", -- 0x1E68
		x"30",x"04",x"3E",x"04",x"18",x"06",x"FE",x"0A", -- 0x1E70
		x"38",x"02",x"3E",x"0A",x"3D",x"E6",x"0F",x"DD", -- 0x1E78
		x"77",x"29",x"CD",x"05",x"58",x"5E",x"FD",x"73", -- 0x1E80
		x"09",x"FD",x"72",x"0A",x"DD",x"7E",x"07",x"FD", -- 0x1E88
		x"77",x"0F",x"DD",x"7E",x"06",x"FD",x"77",x"0E", -- 0x1E90
		x"16",x"02",x"C6",x"05",x"FE",x"7C",x"38",x"07", -- 0x1E98
		x"15",x"FE",x"80",x"30",x"02",x"16",x"03",x"7B", -- 0x1EA0
		x"06",x"01",x"1E",x"02",x"FE",x"06",x"38",x"05", -- 0x1EA8
		x"04",x"FE",x"08",x"38",x"0A",x"A0",x"20",x"01", -- 0x1EB0
		x"1D",x"7B",x"BA",x"28",x"02",x"16",x"03",x"CD", -- 0x1EB8
		x"51",x"0C",x"D8",x"CD",x"31",x"5F",x"FD",x"77", -- 0x1EC0
		x"0B",x"FD",x"4E",x"09",x"79",x"E6",x"FE",x"FE", -- 0x1EC8
		x"06",x"16",x"00",x"28",x"01",x"14",x"3A",x"04", -- 0x1ED0
		x"C0",x"E6",x"60",x"21",x"00",x"78",x"20",x"03", -- 0x1ED8
		x"21",x"40",x"78",x"CB",x"01",x"CB",x"01",x"06", -- 0x1EE0
		x"00",x"09",x"3A",x"0C",x"E0",x"07",x"07",x"E6", -- 0x1EE8
		x"1F",x"5F",x"7E",x"83",x"FD",x"77",x"07",x"23", -- 0x1EF0
		x"7E",x"FD",x"77",x"08",x"23",x"3A",x"F0",x"E0", -- 0x1EF8
		x"2F",x"32",x"F0",x"E0",x"83",x"E6",x"1F",x"5F", -- 0x1F00
		x"7E",x"CB",x"42",x"28",x"01",x"83",x"FD",x"77", -- 0x1F08
		x"05",x"23",x"7E",x"FD",x"77",x"06",x"FD",x"36", -- 0x1F10
		x"0C",x"BB",x"FD",x"36",x"0D",x"0E",x"FD",x"4E", -- 0x1F18
		x"09",x"21",x"37",x"5F",x"09",x"7E",x"FD",x"77", -- 0x1F20
		x"09",x"AF",x"FD",x"77",x"03",x"FD",x"77",x"04", -- 0x1F28
		x"C9",x"7D",x"E6",x"1F",x"07",x"07",x"C9",x"02", -- 0x1F30
		x"03",x"00",x"01",x"00",x"01",x"02",x"00",x"02", -- 0x1F38
		x"02",x"03",x"03",x"00",x"00",x"01",x"01",x"06", -- 0x1F40
		x"09",x"00",x"08",x"04",x"0C",x"02",x"0D",x"07", -- 0x1F48
		x"0F",x"03",x"0E",x"05",x"0A",x"01",x"0B",x"2A", -- 0x1F50
		x"0E",x"E1",x"7D",x"DD",x"BE",x"06",x"30",x"14", -- 0x1F58
		x"C6",x"1F",x"DD",x"BE",x"06",x"38",x"0D",x"1E", -- 0x1F60
		x"07",x"7C",x"C6",x"08",x"DD",x"BE",x"07",x"30", -- 0x1F68
		x"44",x"1D",x"18",x"41",x"7C",x"DD",x"BE",x"07", -- 0x1F70
		x"30",x"14",x"C6",x"0F",x"DD",x"BE",x"07",x"38", -- 0x1F78
		x"0D",x"1E",x"05",x"7D",x"C6",x"10",x"DD",x"BE", -- 0x1F80
		x"06",x"38",x"2A",x"1D",x"18",x"27",x"1E",x"02", -- 0x1F88
		x"7D",x"DD",x"96",x"06",x"30",x"03",x"1C",x"ED", -- 0x1F90
		x"44",x"6F",x"E6",x"F0",x"4F",x"7C",x"DD",x"96", -- 0x1F98
		x"07",x"30",x"04",x"1D",x"1D",x"ED",x"44",x"67", -- 0x1FA0
		x"E6",x"F0",x"B9",x"28",x"08",x"CB",x"03",x"CB", -- 0x1FA8
		x"DB",x"B9",x"38",x"01",x"1C",x"3A",x"6A",x"E1", -- 0x1FB0
		x"4F",x"C9",x"CD",x"79",x"60",x"DA",x"0C",x"60", -- 0x1FB8
		x"DD",x"CB",x"02",x"DE",x"DD",x"CB",x"02",x"A6", -- 0x1FC0
		x"0E",x"07",x"CD",x"78",x"11",x"AF",x"67",x"6F", -- 0x1FC8
		x"22",x"7A",x"E0",x"22",x"7C",x"E0",x"DD",x"36", -- 0x1FD0
		x"0C",x"B0",x"DD",x"36",x"0D",x"4E",x"3E",x"01", -- 0x1FD8
		x"32",x"7C",x"E0",x"21",x"7F",x"E0",x"CD",x"D1", -- 0x1FE0
		x"12",x"CD",x"55",x"2D",x"CD",x"E8",x"2A",x"DD", -- 0x1FE8
		x"36",x"13",x"30",x"DD",x"34",x"03",x"DD",x"7E", -- 0x1FF0
		x"02",x"E6",x"07",x"CD",x"F7",x"66",x"B7",x"60", -- 0x1FF8
		x"A5",x"60",x"78",x"61",x"5C",x"61",x"96",x"60", -- 0x2000
		x"B0",x"60",x"77",x"61",x"DD",x"7E",x"15",x"B7", -- 0x2008
		x"28",x"0F",x"DD",x"35",x"15",x"20",x"0A",x"DD", -- 0x2010
		x"7E",x"16",x"DD",x"77",x"0C",x"DD",x"36",x"0D", -- 0x2018
		x"0E",x"DD",x"CB",x"0D",x"66",x"CA",x"3D",x"60", -- 0x2020
		x"DD",x"7E",x"0F",x"FE",x"F1",x"D2",x"3D",x"60", -- 0x2028
		x"DD",x"CB",x"02",x"DE",x"CD",x"CB",x"66",x"3E", -- 0x2030
		x"01",x"32",x"EA",x"E7",x"C9",x"DD",x"CB",x"02", -- 0x2038
		x"66",x"CA",x"DE",x"61",x"DD",x"6E",x"10",x"DD", -- 0x2040
		x"66",x"11",x"4E",x"23",x"7E",x"DD",x"CB",x"02", -- 0x2048
		x"6E",x"C4",x"90",x"39",x"47",x"CD",x"FB",x"3A", -- 0x2050
		x"D8",x"DD",x"35",x"16",x"C2",x"E8",x"2A",x"23", -- 0x2058
		x"7E",x"B7",x"28",x"0E",x"DD",x"77",x"16",x"23", -- 0x2060
		x"23",x"DD",x"75",x"10",x"DD",x"74",x"11",x"C3", -- 0x2068
		x"E8",x"2A",x"DD",x"36",x"16",x"FF",x"C3",x"E8", -- 0x2070
		x"2A",x"2A",x"0E",x"E1",x"DD",x"7E",x"0E",x"5F", -- 0x2078
		x"C6",x"0F",x"BD",x"D8",x"7D",x"C6",x"1F",x"BB", -- 0x2080
		x"D8",x"DD",x"7E",x"0F",x"57",x"C6",x"0F",x"BC", -- 0x2088
		x"D8",x"7C",x"C6",x"0F",x"BA",x"C9",x"DD",x"CB", -- 0x2090
		x"02",x"7E",x"CA",x"C5",x"2D",x"3E",x"01",x"32", -- 0x2098
		x"13",x"E1",x"C3",x"C5",x"2D",x"21",x"64",x"E1", -- 0x20A0
		x"CB",x"FE",x"21",x"1F",x"E1",x"CB",x"CE",x"C9", -- 0x20A8
		x"21",x"9B",x"E0",x"34",x"C3",x"67",x"18",x"21", -- 0x20B0
		x"00",x"00",x"22",x"78",x"E0",x"22",x"7A",x"E0", -- 0x20B8
		x"22",x"7C",x"E0",x"22",x"7E",x"E0",x"FD",x"21", -- 0x20C0
		x"00",x"E4",x"06",x"10",x"C5",x"FD",x"7E",x"00", -- 0x20C8
		x"57",x"E6",x"07",x"FE",x"01",x"20",x"47",x"FD", -- 0x20D0
		x"7E",x"03",x"B7",x"28",x"41",x"7A",x"E6",x"C0", -- 0x20D8
		x"FE",x"80",x"30",x"3A",x"CB",x"72",x"FD",x"7E", -- 0x20E0
		x"01",x"20",x"15",x"E6",x"C0",x"07",x"07",x"07", -- 0x20E8
		x"4F",x"06",x"00",x"21",x"4C",x"61",x"09",x"7E", -- 0x20F0
		x"23",x"66",x"6F",x"0E",x"07",x"09",x"18",x"0A", -- 0x20F8
		x"FD",x"7E",x"13",x"FE",x"05",x"30",x"17",x"21", -- 0x2100
		x"5B",x"61",x"FD",x"CB",x"00",x"CE",x"11",x"7F", -- 0x2108
		x"E0",x"06",x"08",x"CD",x"FA",x"01",x"21",x"70", -- 0x2110
		x"E1",x"7E",x"B7",x"28",x"01",x"35",x"01",x"30", -- 0x2118
		x"00",x"FD",x"09",x"C1",x"10",x"A6",x"21",x"7F", -- 0x2120
		x"E0",x"CD",x"D1",x"12",x"CD",x"55",x"2D",x"FD", -- 0x2128
		x"21",x"00",x"E3",x"06",x"0F",x"11",x"10",x"00", -- 0x2130
		x"FD",x"7E",x"00",x"CB",x"47",x"28",x"08",x"CB", -- 0x2138
		x"4F",x"20",x"04",x"FD",x"CB",x"00",x"D6",x"FD", -- 0x2140
		x"19",x"10",x"ED",x"C9",x"54",x"38",x"5C",x"38", -- 0x2148
		x"7C",x"38",x"32",x"38",x"00",x"00",x"00",x"00", -- 0x2150
		x"02",x"00",x"00",x"00",x"21",x"0F",x"3C",x"22", -- 0x2158
		x"A2",x"E9",x"21",x"C2",x"E0",x"F3",x"CB",x"4E", -- 0x2160
		x"20",x"08",x"36",x"02",x"FB",x"DD",x"36",x"14", -- 0x2168
		x"01",x"C9",x"FB",x"DD",x"36",x"14",x"00",x"C9", -- 0x2170
		x"AF",x"32",x"20",x"E1",x"3E",x"40",x"32",x"30", -- 0x2178
		x"E1",x"3E",x"03",x"32",x"18",x"E1",x"21",x"1F", -- 0x2180
		x"E1",x"CB",x"C6",x"C9",x"CD",x"94",x"61",x"DD", -- 0x2188
		x"36",x"00",x"00",x"C9",x"AF",x"DD",x"77",x"0D", -- 0x2190
		x"DD",x"77",x"0E",x"CD",x"E8",x"2A",x"C3",x"02", -- 0x2198
		x"67",x"DD",x"7E",x"02",x"E6",x"07",x"FE",x"03", -- 0x21A0
		x"28",x"07",x"DD",x"35",x"13",x"C0",x"C3",x"8C", -- 0x21A8
		x"61",x"DD",x"7E",x"13",x"B7",x"28",x"15",x"DD", -- 0x21B0
		x"35",x"13",x"28",x"07",x"DD",x"7E",x"14",x"B7", -- 0x21B8
		x"C8",x"18",x"09",x"CD",x"94",x"61",x"DD",x"7E", -- 0x21C0
		x"14",x"B7",x"28",x"0E",x"21",x"A3",x"E9",x"35", -- 0x21C8
		x"C0",x"36",x"3C",x"2B",x"35",x"C0",x"AF",x"32", -- 0x21D0
		x"C2",x"E0",x"DD",x"77",x"00",x"C9",x"3A",x"C7", -- 0x21D8
		x"EB",x"CB",x"4F",x"28",x"21",x"DD",x"7E",x"0D", -- 0x21E0
		x"E6",x"10",x"28",x"02",x"3E",x"01",x"67",x"DD", -- 0x21E8
		x"6E",x"0F",x"2B",x"DD",x"75",x"0F",x"7C",x"E6", -- 0x21F0
		x"01",x"28",x"07",x"DD",x"CB",x"0D",x"E6",x"C3", -- 0x21F8
		x"E8",x"2A",x"DD",x"CB",x"0D",x"A6",x"C3",x"E8", -- 0x2200
		x"2A",x"DD",x"CB",x"0D",x"66",x"DD",x"6E",x"0F", -- 0x2208
		x"26",x"00",x"C8",x"24",x"C9",x"DD",x"E5",x"D1", -- 0x2210
		x"7A",x"E6",x"01",x"B3",x"07",x"07",x"07",x"E6", -- 0x2218
		x"0F",x"21",x"E0",x"E0",x"B5",x"6F",x"C9",x"CB", -- 0x2220
		x"57",x"C2",x"83",x"63",x"57",x"E6",x"C0",x"FE", -- 0x2228
		x"40",x"28",x"1F",x"DD",x"7E",x"01",x"E6",x"C0", -- 0x2230
		x"FE",x"C0",x"28",x"16",x"DD",x"7E",x"08",x"E6", -- 0x2238
		x"C0",x"FE",x"80",x"20",x"0D",x"DD",x"6E",x"22", -- 0x2240
		x"DD",x"66",x"23",x"E5",x"FD",x"E1",x"FD",x"CB", -- 0x2248
		x"02",x"A6",x"DD",x"CB",x"00",x"E6",x"DD",x"CB", -- 0x2250
		x"00",x"D6",x"DD",x"36",x"1C",x"00",x"7A",x"E6", -- 0x2258
		x"C0",x"FE",x"40",x"CA",x"F2",x"62",x"FE",x"C0", -- 0x2260
		x"CA",x"44",x"63",x"DD",x"7E",x"01",x"E6",x"C0", -- 0x2268
		x"FE",x"C0",x"CA",x"B1",x"62",x"3A",x"03",x"E1", -- 0x2270
		x"FE",x"01",x"38",x"11",x"21",x"04",x"E1",x"35", -- 0x2278
		x"20",x"0B",x"36",x"C8",x"21",x"09",x"E1",x"34", -- 0x2280
		x"21",x"07",x"E1",x"CB",x"C6",x"DD",x"36",x"0C", -- 0x2288
		x"D8",x"DD",x"7E",x"0D",x"E6",x"10",x"F6",x"0E", -- 0x2290
		x"DD",x"77",x"0D",x"CD",x"E8",x"2A",x"DD",x"36", -- 0x2298
		x"13",x"02",x"3A",x"A5",x"E0",x"0F",x"DA",x"23", -- 0x22A0
		x"2F",x"0E",x"04",x"CD",x"78",x"11",x"C3",x"23", -- 0x22A8
		x"2F",x"3E",x"E8",x"DD",x"77",x"2C",x"C6",x"02", -- 0x22B0
		x"DD",x"77",x"0C",x"DD",x"7E",x"2E",x"DD",x"77", -- 0x22B8
		x"0E",x"DD",x"7E",x"1A",x"C6",x"26",x"57",x"DD", -- 0x22C0
		x"7E",x"2D",x"E6",x"50",x"B2",x"DD",x"77",x"2D", -- 0x22C8
		x"DD",x"7E",x"0D",x"E6",x"50",x"B2",x"DD",x"77", -- 0x22D0
		x"0D",x"CD",x"E8",x"2A",x"CD",x"D9",x"4F",x"DD", -- 0x22D8
		x"36",x"13",x"03",x"3A",x"A5",x"E0",x"0F",x"DA", -- 0x22E0
		x"23",x"2F",x"0E",x"04",x"CD",x"78",x"11",x"C3", -- 0x22E8
		x"23",x"2F",x"DD",x"CB",x"01",x"76",x"C2",x"65", -- 0x22F0
		x"63",x"DD",x"7E",x"1A",x"C6",x"06",x"4F",x"06", -- 0x22F8
		x"F0",x"DD",x"7E",x"0D",x"A0",x"B1",x"DD",x"77", -- 0x2300
		x"0D",x"3A",x"13",x"EC",x"A0",x"B1",x"32",x"13", -- 0x2308
		x"EC",x"3A",x"18",x"EC",x"A0",x"B1",x"32",x"18", -- 0x2310
		x"EC",x"3A",x"1D",x"EC",x"A0",x"B1",x"32",x"1D", -- 0x2318
		x"EC",x"3E",x"07",x"32",x"02",x"EC",x"CD",x"7B", -- 0x2320
		x"53",x"CD",x"1A",x"54",x"DD",x"36",x"13",x"05", -- 0x2328
		x"3A",x"A5",x"E0",x"0F",x"DA",x"AE",x"65",x"3E", -- 0x2330
		x"0B",x"CD",x"78",x"11",x"0E",x"02",x"CD",x"78", -- 0x2338
		x"11",x"C3",x"AE",x"65",x"DD",x"36",x"13",x"02", -- 0x2340
		x"21",x"3E",x"A1",x"DD",x"75",x"10",x"DD",x"74", -- 0x2348
		x"11",x"7E",x"DD",x"77",x"14",x"DD",x"7E",x"00", -- 0x2350
		x"E6",x"C1",x"F6",x"10",x"DD",x"77",x"00",x"DD", -- 0x2358
		x"34",x"03",x"C3",x"23",x"2F",x"21",x"D0",x"EB", -- 0x2360
		x"CB",x"E6",x"3E",x"03",x"32",x"D4",x"E9",x"3E", -- 0x2368
		x"02",x"32",x"F8",x"E9",x"21",x"56",x"7F",x"22", -- 0x2370
		x"FE",x"E9",x"CD",x"68",x"66",x"CD",x"A6",x"5C", -- 0x2378
		x"C3",x"99",x"30",x"CB",x"77",x"C2",x"3F",x"65", -- 0x2380
		x"DD",x"7E",x"01",x"2F",x"E6",x"C0",x"CA",x"BE", -- 0x2388
		x"63",x"DD",x"35",x"13",x"C2",x"23",x"2F",x"DD", -- 0x2390
		x"7E",x"1C",x"3C",x"FE",x"06",x"D2",x"4C",x"64", -- 0x2398
		x"DD",x"77",x"1C",x"21",x"B8",x"63",x"4F",x"06", -- 0x23A0
		x"00",x"09",x"7E",x"DD",x"77",x"0C",x"CD",x"E8", -- 0x23A8
		x"2A",x"DD",x"36",x"13",x"04",x"C3",x"23",x"2F", -- 0x23B0
		x"D8",x"D9",x"DA",x"DB",x"DC",x"DD",x"DD",x"35", -- 0x23B8
		x"13",x"C2",x"23",x"2F",x"DD",x"7E",x"1C",x"3C", -- 0x23C0
		x"FE",x"0A",x"D2",x"E8",x"63",x"DD",x"77",x"1C", -- 0x23C8
		x"CD",x"2E",x"64",x"DD",x"77",x"2C",x"23",x"7E", -- 0x23D0
		x"DD",x"77",x"0C",x"CD",x"E8",x"2A",x"CD",x"D9", -- 0x23D8
		x"4F",x"DD",x"36",x"13",x"05",x"C3",x"23",x"2F", -- 0x23E0
		x"FE",x"0B",x"30",x"3D",x"DD",x"77",x"1C",x"DD", -- 0x23E8
		x"7E",x"1D",x"B7",x"01",x"B1",x"B0",x"28",x"03", -- 0x23F0
		x"01",x"D7",x"B0",x"DD",x"70",x"0C",x"DD",x"71", -- 0x23F8
		x"2C",x"DD",x"7E",x"0D",x"E6",x"10",x"F6",x"0E", -- 0x2400
		x"DD",x"77",x"0D",x"DD",x"77",x"2D",x"DD",x"7E", -- 0x2408
		x"0E",x"C6",x"10",x"DD",x"77",x"2E",x"DD",x"7E", -- 0x2410
		x"0F",x"DD",x"77",x"2F",x"CD",x"E8",x"2A",x"CD", -- 0x2418
		x"D9",x"4F",x"DD",x"36",x"13",x"14",x"C3",x"23", -- 0x2420
		x"2F",x"CD",x"DD",x"66",x"18",x"2E",x"21",x"38", -- 0x2428
		x"64",x"07",x"4F",x"06",x"00",x"09",x"7E",x"C9", -- 0x2430
		x"E8",x"EA",x"EC",x"EE",x"E8",x"EA",x"F0",x"F2", -- 0x2438
		x"E8",x"EA",x"EC",x"EE",x"F0",x"F2",x"F4",x"F6", -- 0x2440
		x"F8",x"FA",x"FC",x"FE",x"DD",x"7E",x"08",x"E6", -- 0x2448
		x"E0",x"20",x"0F",x"DD",x"CB",x"01",x"6E",x"28", -- 0x2450
		x"03",x"CD",x"FD",x"64",x"CD",x"CB",x"66",x"C3", -- 0x2458
		x"23",x"2F",x"DD",x"6E",x"1E",x"DD",x"66",x"1F", -- 0x2460
		x"35",x"23",x"C2",x"F3",x"64",x"35",x"01",x"4E", -- 0x2468
		x"B0",x"21",x"39",x"65",x"FE",x"60",x"28",x"05", -- 0x2470
		x"21",x"3E",x"65",x"06",x"B2",x"DD",x"70",x"0C", -- 0x2478
		x"DD",x"71",x"0D",x"CD",x"D1",x"12",x"CD",x"55", -- 0x2480
		x"2D",x"AF",x"47",x"57",x"DD",x"7E",x"08",x"E6", -- 0x2488
		x"E0",x"FE",x"60",x"DD",x"7E",x"02",x"20",x"08", -- 0x2490
		x"E6",x"0F",x"FE",x"05",x"28",x"29",x"18",x"25", -- 0x2498
		x"E6",x"0F",x"FE",x"04",x"20",x"04",x"3E",x"84", -- 0x24A0
		x"18",x"1D",x"FE",x"02",x"20",x"0A",x"3A",x"1F", -- 0x24A8
		x"E1",x"0F",x"38",x"11",x"3E",x"02",x"18",x"0F", -- 0x24B0
		x"FE",x"01",x"20",x"0B",x"3A",x"1F",x"E1",x"CB", -- 0x24B8
		x"4F",x"3E",x"01",x"28",x"02",x"3E",x"06",x"DD", -- 0x24C0
		x"77",x"02",x"E6",x"07",x"06",x"00",x"4F",x"21", -- 0x24C8
		x"2B",x"65",x"09",x"7E",x"DD",x"77",x"16",x"AF", -- 0x24D0
		x"32",x"EA",x"E7",x"DD",x"77",x"17",x"DD",x"77", -- 0x24D8
		x"03",x"DD",x"36",x"15",x"14",x"DD",x"36",x"13", -- 0x24E0
		x"D2",x"DD",x"36",x"00",x"81",x"CD",x"E8",x"2A", -- 0x24E8
		x"C3",x"23",x"2F",x"35",x"C2",x"5C",x"64",x"CD", -- 0x24F0
		x"25",x"65",x"C3",x"23",x"2F",x"21",x"1E",x"E1", -- 0x24F8
		x"7E",x"B7",x"28",x"01",x"35",x"7E",x"47",x"21", -- 0x2500
		x"1D",x"E1",x"F3",x"BE",x"30",x"0D",x"96",x"ED", -- 0x2508
		x"44",x"32",x"1B",x"E1",x"21",x"1E",x"E1",x"86", -- 0x2510
		x"77",x"FB",x"C9",x"7E",x"B7",x"20",x"FA",x"AF", -- 0x2518
		x"32",x"1E",x"E1",x"18",x"F4",x"CD",x"37",x"60", -- 0x2520
		x"C3",x"CB",x"66",x"0F",x"3F",x"2F",x"3B",x"1F", -- 0x2528
		x"C6",x"C7",x"00",x"00",x"00",x"00",x"01",x"00", -- 0x2530
		x"00",x"00",x"00",x"00",x"05",x"00",x"00",x"DD", -- 0x2538
		x"CB",x"01",x"76",x"C2",x"BA",x"65",x"DD",x"35", -- 0x2540
		x"13",x"C2",x"AE",x"65",x"DD",x"7E",x"1C",x"3C", -- 0x2548
		x"FE",x"09",x"30",x"1A",x"DD",x"77",x"1C",x"4F", -- 0x2550
		x"06",x"00",x"21",x"B1",x"65",x"09",x"7E",x"32", -- 0x2558
		x"02",x"EC",x"CD",x"7B",x"53",x"CD",x"1A",x"54", -- 0x2560
		x"DD",x"36",x"13",x"07",x"18",x"40",x"3A",x"13", -- 0x2568
		x"EC",x"E6",x"0F",x"D6",x"06",x"07",x"4F",x"3A", -- 0x2570
		x"13",x"EC",x"E6",x"F0",x"B1",x"32",x"13",x"EC", -- 0x2578
		x"3A",x"18",x"EC",x"E6",x"F0",x"B1",x"32",x"18", -- 0x2580
		x"EC",x"3E",x"02",x"32",x"02",x"EC",x"CD",x"7B", -- 0x2588
		x"53",x"CD",x"1A",x"54",x"DD",x"7E",x"00",x"E6", -- 0x2590
		x"F9",x"F6",x"18",x"DD",x"77",x"00",x"DD",x"36", -- 0x2598
		x"15",x"04",x"DD",x"36",x"16",x"08",x"DD",x"36", -- 0x25A0
		x"13",x"05",x"DD",x"36",x"03",x"02",x"C3",x"23", -- 0x25A8
		x"2F",x"07",x"08",x"09",x"0A",x"08",x"09",x"0A", -- 0x25B0
		x"0B",x"0C",x"CD",x"A6",x"5C",x"CD",x"60",x"66", -- 0x25B8
		x"D2",x"99",x"30",x"21",x"00",x"E3",x"01",x"00", -- 0x25C0
		x"0F",x"11",x"10",x"00",x"71",x"19",x"10",x"FC", -- 0x25C8
		x"21",x"11",x"EB",x"06",x"1C",x"71",x"23",x"71", -- 0x25D0
		x"23",x"23",x"23",x"10",x"F8",x"21",x"A4",x"EB", -- 0x25D8
		x"06",x"1C",x"71",x"23",x"10",x"FC",x"11",x"50", -- 0x25E0
		x"EB",x"21",x"50",x"66",x"01",x"0C",x"00",x"ED", -- 0x25E8
		x"B0",x"11",x"70",x"EB",x"21",x"50",x"66",x"01", -- 0x25F0
		x"0C",x"00",x"ED",x"B0",x"3A",x"03",x"E1",x"E6", -- 0x25F8
		x"18",x"0F",x"0F",x"0F",x"4F",x"06",x"00",x"21", -- 0x2600
		x"5C",x"66",x"09",x"7E",x"32",x"50",x"EB",x"32", -- 0x2608
		x"70",x"EB",x"DD",x"7E",x"0F",x"C6",x"40",x"32", -- 0x2610
		x"53",x"EB",x"32",x"57",x"EB",x"32",x"5B",x"EB", -- 0x2618
		x"32",x"73",x"EB",x"32",x"77",x"EB",x"32",x"7B", -- 0x2620
		x"EB",x"DD",x"7E",x"00",x"E6",x"F9",x"F6",x"10", -- 0x2628
		x"DD",x"77",x"00",x"DD",x"36",x"14",x"3C",x"DD", -- 0x2630
		x"36",x"13",x"00",x"DD",x"36",x"03",x"02",x"AF", -- 0x2638
		x"32",x"B4",x"E7",x"0E",x"0B",x"CD",x"78",x"11", -- 0x2640
		x"0E",x"15",x"CD",x"78",x"11",x"C3",x"99",x"30", -- 0x2648
		x"47",x"0E",x"68",x"00",x"B1",x"0E",x"78",x"00", -- 0x2650
		x"B4",x"0E",x"87",x"00",x"47",x"4B",x"4F",x"B2", -- 0x2658
		x"21",x"FB",x"E9",x"35",x"C0",x"2A",x"FE",x"E9", -- 0x2660
		x"7E",x"B7",x"CA",x"BF",x"66",x"47",x"23",x"7E", -- 0x2668
		x"32",x"FB",x"E9",x"23",x"DD",x"7E",x"0F",x"86", -- 0x2670
		x"DD",x"77",x"07",x"23",x"DD",x"7E",x"0E",x"86", -- 0x2678
		x"DD",x"77",x"06",x"23",x"CD",x"11",x"67",x"38", -- 0x2680
		x"29",x"D9",x"CD",x"51",x"0C",x"7D",x"D9",x"38", -- 0x2688
		x"28",x"CD",x"32",x"5F",x"FD",x"77",x"0B",x"3A", -- 0x2690
		x"F0",x"E3",x"3C",x"32",x"F0",x"E3",x"DD",x"7E", -- 0x2698
		x"07",x"FD",x"77",x"0F",x"DD",x"7E",x"06",x"FD", -- 0x26A0
		x"77",x"0E",x"FD",x"36",x"0D",x"0E",x"FD",x"36", -- 0x26A8
		x"00",x"09",x"10",x"C0",x"22",x"FE",x"E9",x"B7", -- 0x26B0
		x"C9",x"FD",x"36",x"00",x"00",x"18",x"F3",x"21", -- 0x26B8
		x"D4",x"E9",x"35",x"21",x"56",x"7F",x"C2",x"68", -- 0x26C0
		x"66",x"37",x"C9",x"AF",x"DD",x"77",x"0D",x"DD", -- 0x26C8
		x"77",x"0E",x"CD",x"E8",x"2A",x"CD",x"02",x"67", -- 0x26D0
		x"DD",x"36",x"00",x"00",x"C9",x"AF",x"DD",x"77", -- 0x26D8
		x"2D",x"DD",x"77",x"2E",x"DD",x"E5",x"E1",x"01", -- 0x26E0
		x"2B",x"00",x"09",x"CD",x"EF",x"2A",x"DD",x"7E", -- 0x26E8
		x"2B",x"C3",x"05",x"67",x"DD",x"7E",x"03",x"07", -- 0x26F0
		x"4F",x"06",x"00",x"E1",x"09",x"7E",x"23",x"66", -- 0x26F8
		x"6F",x"E9",x"DD",x"7E",x"0B",x"21",x"A0",x"EB", -- 0x2700
		x"0F",x"0F",x"E6",x"1F",x"B5",x"6F",x"CB",x"BE", -- 0x2708
		x"C9",x"B7",x"D9",x"FD",x"21",x"00",x"E3",x"06", -- 0x2710
		x"0F",x"11",x"10",x"00",x"FD",x"7E",x"00",x"E6", -- 0x2718
		x"03",x"20",x"06",x"FD",x"CB",x"00",x"CE",x"D9", -- 0x2720
		x"C9",x"FD",x"19",x"10",x"EF",x"D9",x"37",x"C9", -- 0x2728
		x"3E",x"01",x"32",x"A5",x"E0",x"3A",x"03",x"E1", -- 0x2730
		x"32",x"06",x"E1",x"3E",x"09",x"EF",x"3E",x"0E", -- 0x2738
		x"EF",x"21",x"00",x"E1",x"CB",x"AE",x"3A",x"00", -- 0x2740
		x"E0",x"07",x"38",x"0B",x"3E",x"0D",x"EF",x"21", -- 0x2748
		x"96",x"A4",x"CD",x"22",x"02",x"18",x"0B",x"21", -- 0x2750
		x"08",x"D0",x"01",x"10",x"1C",x"16",x"30",x"CD", -- 0x2758
		x"53",x"02",x"21",x"FF",x"FF",x"22",x"72",x"E1", -- 0x2760
		x"22",x"72",x"E1",x"3E",x"01",x"32",x"76",x"E1", -- 0x2768
		x"0E",x"00",x"CD",x"78",x"11",x"0E",x"0F",x"CD", -- 0x2770
		x"78",x"11",x"0E",x"0B",x"CD",x"78",x"11",x"0E", -- 0x2778
		x"10",x"CD",x"78",x"11",x"0E",x"02",x"CD",x"78", -- 0x2780
		x"11",x"AF",x"67",x"6F",x"22",x"05",x"EB",x"22", -- 0x2788
		x"09",x"EB",x"22",x"0D",x"EB",x"32",x"60",x"E2", -- 0x2790
		x"32",x"70",x"E2",x"32",x"80",x"E2",x"3A",x"B4", -- 0x2798
		x"E7",x"B7",x"20",x"1F",x"21",x"48",x"EB",x"11", -- 0x27A0
		x"49",x"EB",x"01",x"17",x"00",x"36",x"00",x"ED", -- 0x27A8
		x"B0",x"21",x"68",x"EB",x"11",x"69",x"EB",x"01", -- 0x27B0
		x"17",x"00",x"36",x"00",x"ED",x"B0",x"06",x"02", -- 0x27B8
		x"DF",x"18",x"14",x"3A",x"A9",x"E0",x"B7",x"28", -- 0x27C0
		x"0E",x"3A",x"A6",x"E9",x"CB",x"4F",x"28",x"07", -- 0x27C8
		x"AF",x"32",x"20",x"E1",x"32",x"30",x"E1",x"21", -- 0x27D0
		x"0C",x"E1",x"11",x"00",x"EB",x"01",x"04",x"00", -- 0x27D8
		x"ED",x"B0",x"21",x"0C",x"E1",x"01",x"04",x"00", -- 0x27E0
		x"ED",x"B0",x"3A",x"0F",x"E1",x"D6",x"08",x"32", -- 0x27E8
		x"03",x"EB",x"C6",x"10",x"32",x"07",x"EB",x"3A", -- 0x27F0
		x"20",x"E1",x"E6",x"82",x"FE",x"80",x"CC",x"E6", -- 0x27F8
		x"68",x"3A",x"30",x"E1",x"E6",x"82",x"FE",x"80", -- 0x2800
		x"CC",x"E0",x"68",x"3E",x"0E",x"32",x"2D",x"E1", -- 0x2808
		x"32",x"3D",x"E1",x"21",x"20",x"E1",x"CB",x"D6", -- 0x2810
		x"21",x"30",x"E1",x"CB",x"D6",x"21",x"84",x"78", -- 0x2818
		x"FD",x"21",x"87",x"87",x"7E",x"B7",x"28",x"44", -- 0x2820
		x"DD",x"21",x"20",x"E1",x"DD",x"7E",x"00",x"2F", -- 0x2828
		x"E6",x"82",x"20",x"0B",x"FD",x"7E",x"01",x"DD", -- 0x2830
		x"77",x"0C",x"E5",x"CD",x"E8",x"2A",x"E1",x"DD", -- 0x2838
		x"7E",x"10",x"2F",x"E6",x"82",x"20",x"12",x"FD", -- 0x2840
		x"7E",x"01",x"DD",x"77",x"1C",x"E5",x"DD",x"E5", -- 0x2848
		x"E1",x"01",x"1B",x"00",x"09",x"CD",x"EF",x"2A", -- 0x2850
		x"E1",x"FD",x"23",x"FD",x"23",x"11",x"00",x"EB", -- 0x2858
		x"ED",x"A0",x"11",x"04",x"EB",x"ED",x"A0",x"46", -- 0x2860
		x"DF",x"23",x"18",x"B8",x"21",x"00",x"00",x"22", -- 0x2868
		x"0C",x"E1",x"22",x"0E",x"E1",x"22",x"04",x"EB", -- 0x2870
		x"22",x"06",x"EB",x"CD",x"3A",x"29",x"DD",x"21", -- 0x2878
		x"20",x"E1",x"AF",x"DD",x"77",x"0D",x"DD",x"77", -- 0x2880
		x"0E",x"DD",x"77",x"1D",x"DD",x"77",x"1E",x"DD", -- 0x2888
		x"CB",x"00",x"7E",x"C4",x"E8",x"2A",x"DD",x"36", -- 0x2890
		x"00",x"00",x"DD",x"21",x"30",x"E1",x"DD",x"CB", -- 0x2898
		x"00",x"7E",x"C4",x"E8",x"2A",x"AF",x"DD",x"77", -- 0x28A0
		x"00",x"3E",x"02",x"EF",x"3C",x"EF",x"0E",x"03", -- 0x28A8
		x"C5",x"06",x"1E",x"DF",x"C1",x"0D",x"20",x"F8", -- 0x28B0
		x"0E",x"00",x"CD",x"78",x"11",x"AF",x"32",x"1F", -- 0x28B8
		x"E1",x"32",x"64",x"E1",x"32",x"07",x"EC",x"3A", -- 0x28C0
		x"00",x"E0",x"07",x"38",x"2C",x"06",x"40",x"DF", -- 0x28C8
		x"3E",x"01",x"EF",x"3E",x"04",x"EF",x"3E",x"05", -- 0x28D0
		x"EF",x"AF",x"32",x"C7",x"EB",x"C3",x"8A",x"0F", -- 0x28D8
		x"DD",x"21",x"30",x"E1",x"18",x"04",x"DD",x"21", -- 0x28E0
		x"20",x"E1",x"DD",x"CB",x"00",x"46",x"C8",x"AF", -- 0x28E8
		x"DD",x"77",x"0D",x"DD",x"77",x"0E",x"C3",x"E8", -- 0x28F0
		x"2A",x"3E",x"04",x"EF",x"21",x"01",x"E1",x"7E", -- 0x28F8
		x"FE",x"01",x"20",x"21",x"DD",x"21",x"A0",x"A2", -- 0x2900
		x"CD",x"CC",x"2C",x"21",x"45",x"A5",x"CD",x"22", -- 0x2908
		x"02",x"AF",x"32",x"A6",x"E9",x"32",x"C7",x"EB", -- 0x2910
		x"3E",x"05",x"01",x"51",x"6F",x"FF",x"0E",x"16", -- 0x2918
		x"CD",x"78",x"11",x"18",x"05",x"3E",x"01",x"32", -- 0x2920
		x"A6",x"E9",x"06",x"08",x"DF",x"3A",x"A6",x"E9", -- 0x2928
		x"0F",x"30",x"F7",x"AF",x"32",x"C7",x"EB",x"21", -- 0x2930
		x"01",x"E1",x"35",x"CA",x"96",x"69",x"CD",x"2F", -- 0x2938
		x"2D",x"3A",x"01",x"E0",x"20",x"01",x"0F",x"0F", -- 0x2940
		x"38",x"02",x"18",x"03",x"CD",x"55",x"69",x"3E", -- 0x2948
		x"01",x"EF",x"C3",x"F2",x"14",x"CD",x"6D",x"6A", -- 0x2950
		x"CD",x"2F",x"2D",x"3E",x"02",x"28",x"01",x"0F", -- 0x2958
		x"32",x"A6",x"E0",x"3A",x"03",x"C0",x"E6",x"08", -- 0x2960
		x"0E",x"00",x"28",x"07",x"CD",x"2F",x"2D",x"28", -- 0x2968
		x"02",x"0E",x"80",x"3A",x"04",x"C0",x"E6",x"10", -- 0x2970
		x"20",x"04",x"79",x"EE",x"80",x"4F",x"F3",x"3A", -- 0x2978
		x"D4",x"E0",x"E6",x"7F",x"B1",x"32",x"D4",x"E0", -- 0x2980
		x"FB",x"C9",x"06",x"08",x"AF",x"BE",x"20",x"04", -- 0x2988
		x"23",x"10",x"FA",x"C9",x"37",x"C9",x"CD",x"22", -- 0x2990
		x"12",x"CD",x"E7",x"2C",x"CD",x"2F",x"2D",x"3A", -- 0x2998
		x"01",x"E0",x"20",x"04",x"E6",x"FE",x"18",x"02", -- 0x29A0
		x"E6",x"FD",x"32",x"01",x"E0",x"21",x"40",x"E0", -- 0x29A8
		x"11",x"9C",x"E9",x"CD",x"08",x"6B",x"21",x"00", -- 0x29B0
		x"E1",x"CB",x"BE",x"CD",x"2F",x"2D",x"11",x"48", -- 0x29B8
		x"E0",x"28",x"03",x"11",x"50",x"E0",x"21",x"40", -- 0x29C0
		x"E0",x"06",x"08",x"CD",x"77",x"6B",x"38",x"05", -- 0x29C8
		x"21",x"00",x"E1",x"CB",x"FE",x"06",x"1E",x"DF", -- 0x29D0
		x"0E",x"10",x"CD",x"78",x"11",x"3A",x"01",x"E0", -- 0x29D8
		x"E6",x"03",x"28",x"06",x"CD",x"8B",x"6A",x"C3", -- 0x29E0
		x"4C",x"69",x"21",x"00",x"E0",x"CB",x"D6",x"AF", -- 0x29E8
		x"32",x"9B",x"E9",x"3E",x"02",x"01",x"7F",x"6A", -- 0x29F0
		x"FF",x"06",x"02",x"DF",x"3A",x"9B",x"E9",x"3C", -- 0x29F8
		x"CA",x"56",x"6A",x"2A",x"10",x"E0",x"7D",x"6C", -- 0x2A00
		x"67",x"B5",x"28",x"ED",x"11",x"FE",x"FF",x"19", -- 0x2A08
		x"38",x"11",x"3A",x"00",x"C0",x"E6",x"01",x"20", -- 0x2A10
		x"E0",x"21",x"C4",x"78",x"CD",x"16",x"12",x"3E", -- 0x2A18
		x"01",x"18",x"0F",x"3A",x"00",x"C0",x"E6",x"02", -- 0x2A20
		x"20",x"E8",x"21",x"C6",x"78",x"CD",x"16",x"12", -- 0x2A28
		x"3E",x"83",x"32",x"01",x"E0",x"3E",x"02",x"EF", -- 0x2A30
		x"3C",x"EF",x"21",x"48",x"E0",x"01",x"30",x"00", -- 0x2A38
		x"50",x"CD",x"E2",x"01",x"3E",x"80",x"32",x"00", -- 0x2A40
		x"E0",x"2A",x"04",x"E0",x"23",x"22",x"04",x"E0", -- 0x2A48
		x"CD",x"9C",x"12",x"C3",x"DF",x"14",x"21",x"00", -- 0x2A50
		x"E0",x"7E",x"E6",x"84",x"77",x"3A",x"00",x"E1", -- 0x2A58
		x"E6",x"01",x"C4",x"6D",x"6A",x"0E",x"00",x"CD", -- 0x2A60
		x"78",x"11",x"C3",x"4B",x"13",x"21",x"00",x"E1", -- 0x2A68
		x"11",x"80",x"E1",x"06",x"80",x"4E",x"1A",x"77", -- 0x2A70
		x"79",x"12",x"23",x"13",x"10",x"F7",x"C9",x"CD", -- 0x2A78
		x"8B",x"6A",x"CD",x"6D",x"6A",x"3E",x"FF",x"32", -- 0x2A80
		x"9B",x"E9",x"F7",x"CD",x"A7",x"02",x"CD",x"90", -- 0x2A88
		x"11",x"CD",x"CA",x"11",x"CD",x"9C",x"12",x"CD", -- 0x2A90
		x"4E",x"19",x"21",x"48",x"E0",x"CD",x"2F",x"2D", -- 0x2A98
		x"28",x"03",x"21",x"50",x"E0",x"22",x"97",x"E9", -- 0x2AA0
		x"3A",x"00",x"E1",x"07",x"30",x"07",x"AF",x"32", -- 0x2AA8
		x"92",x"E9",x"C3",x"FC",x"6A",x"11",x"9C",x"E9", -- 0x2AB0
		x"CD",x"08",x"6B",x"3E",x"18",x"32",x"92",x"E9", -- 0x2AB8
		x"CD",x"4C",x"6B",x"23",x"11",x"9C",x"E9",x"CD", -- 0x2AC0
		x"75",x"6B",x"3A",x"92",x"E9",x"30",x"13",x"FE", -- 0x2AC8
		x"18",x"C8",x"3C",x"32",x"92",x"E9",x"FE",x"05", -- 0x2AD0
		x"38",x"22",x"CD",x"1D",x"6B",x"CD",x"7F",x"6B", -- 0x2AD8
		x"18",x"20",x"B7",x"28",x"06",x"3D",x"32",x"92", -- 0x2AE0
		x"E9",x"18",x"D5",x"2A",x"97",x"E9",x"11",x"40", -- 0x2AE8
		x"E0",x"01",x"08",x"00",x"ED",x"B0",x"CD",x"9C", -- 0x2AF0
		x"12",x"CD",x"4E",x"19",x"CD",x"1D",x"6B",x"CD", -- 0x2AF8
		x"85",x"6C",x"21",x"00",x"E0",x"CB",x"86",x"C9", -- 0x2B00
		x"06",x"04",x"7E",x"E6",x"0F",x"07",x"07",x"07", -- 0x2B08
		x"07",x"4F",x"23",x"7E",x"E6",x"0F",x"B1",x"12", -- 0x2B10
		x"23",x"13",x"10",x"EE",x"C9",x"21",x"00",x"E0", -- 0x2B18
		x"CB",x"C6",x"CD",x"E0",x"11",x"3E",x"18",x"CD", -- 0x2B20
		x"4C",x"6B",x"36",x"FE",x"CD",x"57",x"6B",x"23", -- 0x2B28
		x"EB",x"21",x"9C",x"E9",x"0E",x"04",x"ED",x"B0", -- 0x2B30
		x"EB",x"16",x"30",x"0E",x"08",x"CD",x"E2",x"01", -- 0x2B38
		x"3A",x"05",x"E1",x"3C",x"FE",x"63",x"38",x"02", -- 0x2B40
		x"3E",x"63",x"77",x"C9",x"11",x"10",x"00",x"21", -- 0x2B48
		x"00",x"E8",x"BE",x"C8",x"19",x"18",x"FB",x"11", -- 0x2B50
		x"10",x"00",x"3A",x"92",x"E9",x"4F",x"06",x"19", -- 0x2B58
		x"21",x"00",x"E8",x"7E",x"B9",x"38",x"01",x"34", -- 0x2B60
		x"19",x"10",x"F8",x"3E",x"FF",x"CD",x"4C",x"6B", -- 0x2B68
		x"3A",x"92",x"E9",x"77",x"C9",x"06",x"04",x"1A", -- 0x2B70
		x"BE",x"C0",x"23",x"13",x"10",x"F9",x"C9",x"DD", -- 0x2B78
		x"21",x"1A",x"A2",x"CD",x"CC",x"2C",x"CD",x"6C", -- 0x2B80
		x"11",x"21",x"21",x"A5",x"CD",x"22",x"02",x"0E", -- 0x2B88
		x"19",x"CD",x"78",x"11",x"CD",x"0E",x"6F",x"06", -- 0x2B90
		x"05",x"DD",x"21",x"8A",x"D0",x"C5",x"F5",x"CD", -- 0x2B98
		x"4C",x"6B",x"CD",x"BF",x"6B",x"F1",x"3C",x"DD", -- 0x2BA0
		x"2B",x"DD",x"2B",x"C1",x"10",x"EF",x"CD",x"28", -- 0x2BA8
		x"6F",x"11",x"C7",x"78",x"06",x"5A",x"CD",x"34", -- 0x2BB0
		x"6F",x"10",x"FB",x"06",x"01",x"DF",x"C9",x"DD", -- 0x2BB8
		x"E5",x"7E",x"3C",x"0E",x"00",x"FE",x"0A",x"38", -- 0x2BC0
		x"05",x"D6",x"0A",x"0C",x"18",x"F7",x"DD",x"77", -- 0x2BC8
		x"20",x"79",x"B7",x"28",x"03",x"DD",x"77",x"00", -- 0x2BD0
		x"01",x"80",x"00",x"DD",x"09",x"23",x"DD",x"E5", -- 0x2BD8
		x"D1",x"EB",x"CD",x"12",x"6C",x"01",x"20",x"00", -- 0x2BE0
		x"09",x"06",x"08",x"CD",x"EE",x"01",x"CD",x"F4", -- 0x2BE8
		x"6B",x"DD",x"E1",x"C9",x"1A",x"01",x"20",x"00", -- 0x2BF0
		x"09",x"48",x"FE",x"0A",x"38",x"05",x"D6",x"0A", -- 0x2BF8
		x"0C",x"18",x"F7",x"47",x"79",x"B7",x"20",x"02", -- 0x2C00
		x"0E",x"30",x"71",x"78",x"01",x"20",x"00",x"09", -- 0x2C08
		x"77",x"C9",x"0E",x"00",x"06",x"08",x"1A",x"CB", -- 0x2C10
		x"40",x"20",x"04",x"0F",x"0F",x"0F",x"0F",x"E6", -- 0x2C18
		x"0F",x"28",x"04",x"CB",x"C1",x"18",x"0D",x"CB", -- 0x2C20
		x"41",x"20",x"09",x"78",x"FE",x"03",x"3E",x"00", -- 0x2C28
		x"38",x"F1",x"3E",x"30",x"77",x"C5",x"01",x"20", -- 0x2C30
		x"00",x"09",x"C1",x"05",x"CB",x"40",x"20",x"D6", -- 0x2C38
		x"13",x"78",x"B7",x"20",x"D1",x"C9",x"AF",x"32", -- 0x2C40
		x"96",x"E9",x"DD",x"21",x"0B",x"D1",x"06",x"05", -- 0x2C48
		x"C5",x"3A",x"96",x"E9",x"CD",x"4C",x"6B",x"23", -- 0x2C50
		x"EB",x"DD",x"E5",x"E1",x"CD",x"12",x"6C",x"01", -- 0x2C58
		x"20",x"00",x"09",x"06",x"08",x"1A",x"77",x"13", -- 0x2C60
		x"C5",x"01",x"20",x"00",x"09",x"C1",x"10",x"F5", -- 0x2C68
		x"CD",x"F4",x"6B",x"C1",x"DD",x"2B",x"DD",x"2B", -- 0x2C70
		x"21",x"96",x"E9",x"7E",x"B7",x"20",x"02",x"DD", -- 0x2C78
		x"2B",x"34",x"10",x"CC",x"C9",x"DD",x"21",x"ED", -- 0x2C80
		x"A2",x"CD",x"CC",x"2C",x"CD",x"0B",x"6D",x"21", -- 0x2C88
		x"EA",x"A4",x"CD",x"22",x"02",x"21",x"AE",x"D0", -- 0x2C90
		x"01",x"01",x"16",x"16",x"35",x"CD",x"53",x"02", -- 0x2C98
		x"CD",x"46",x"6C",x"3A",x"92",x"E9",x"CD",x"4C", -- 0x2CA0
		x"6B",x"E5",x"DD",x"E1",x"AF",x"32",x"A5",x"E9", -- 0x2CA8
		x"21",x"2B",x"D2",x"3A",x"92",x"E9",x"B7",x"28", -- 0x2CB0
		x"06",x"2B",x"07",x"4F",x"7D",x"91",x"6F",x"22", -- 0x2CB8
		x"90",x"E9",x"01",x"DA",x"6E",x"3E",x"04",x"FF", -- 0x2CC0
		x"01",x"EB",x"6E",x"3E",x"03",x"FF",x"0E",x"17", -- 0x2CC8
		x"CD",x"78",x"11",x"CD",x"3C",x"6D",x"06",x"01", -- 0x2CD0
		x"DF",x"3A",x"A5",x"E9",x"B7",x"28",x"F7",x"0E", -- 0x2CD8
		x"10",x"CD",x"78",x"11",x"3A",x"92",x"E9",x"B7", -- 0x2CE0
		x"28",x"0A",x"0E",x"19",x"CD",x"78",x"11",x"06", -- 0x2CE8
		x"A5",x"DF",x"18",x"08",x"0E",x"18",x"CD",x"78", -- 0x2CF0
		x"11",x"06",x"D5",x"DF",x"06",x"D4",x"DF",x"0E", -- 0x2CF8
		x"10",x"CD",x"78",x"11",x"3E",x"03",x"EF",x"3E", -- 0x2D00
		x"04",x"EF",x"C9",x"21",x"D9",x"D0",x"16",x"0A", -- 0x2D08
		x"06",x"04",x"0E",x"0A",x"E5",x"78",x"3D",x"20", -- 0x2D10
		x"05",x"79",x"FE",x"04",x"38",x"11",x"72",x"14", -- 0x2D18
		x"C5",x"01",x"40",x"00",x"09",x"C1",x"0D",x"20", -- 0x2D20
		x"EC",x"E1",x"2B",x"2B",x"05",x"18",x"E3",x"C1", -- 0x2D28
		x"11",x"20",x"00",x"19",x"19",x"36",x"3B",x"19", -- 0x2D30
		x"19",x"36",x"3D",x"C9",x"21",x"B5",x"00",x"22", -- 0x2D38
		x"00",x"EB",x"21",x"2C",x"C4",x"22",x"02",x"EB", -- 0x2D40
		x"3A",x"92",x"E9",x"CD",x"4C",x"6B",x"E5",x"DD", -- 0x2D48
		x"E1",x"AF",x"32",x"96",x"E9",x"32",x"A0",x"E0", -- 0x2D50
		x"32",x"A3",x"E0",x"32",x"9B",x"E9",x"32",x"A4", -- 0x2D58
		x"E0",x"21",x"03",x"00",x"22",x"94",x"E9",x"3E", -- 0x2D60
		x"1E",x"32",x"93",x"E9",x"CD",x"35",x"2D",x"4F", -- 0x2D68
		x"E6",x"30",x"C2",x"1B",x"6E",x"32",x"A4",x"E0", -- 0x2D70
		x"3A",x"96",x"E9",x"57",x"79",x"E6",x"0F",x"CA", -- 0x2D78
		x"9B",x"6D",x"47",x"3A",x"A0",x"E0",x"B8",x"28", -- 0x2D80
		x"08",x"78",x"32",x"A0",x"E0",x"3E",x"01",x"18", -- 0x2D88
		x"0A",x"3A",x"A3",x"E0",x"3C",x"FE",x"18",x"38", -- 0x2D90
		x"02",x"3E",x"14",x"32",x"A3",x"E0",x"FE",x"01", -- 0x2D98
		x"28",x"07",x"FE",x"14",x"28",x"03",x"7A",x"18", -- 0x2DA0
		x"45",x"79",x"E6",x"0C",x"28",x"1C",x"E6",x"08", -- 0x2DA8
		x"7A",x"28",x"0C",x"FE",x"0A",x"30",x"04",x"C6", -- 0x2DB0
		x"1E",x"18",x"0E",x"D6",x"0A",x"18",x"0A",x"FE", -- 0x2DB8
		x"1E",x"38",x"04",x"D6",x"1E",x"18",x"02",x"C6", -- 0x2DC0
		x"0A",x"57",x"79",x"E6",x"03",x"7A",x"28",x"1E", -- 0x2DC8
		x"79",x"E6",x"02",x"7A",x"28",x"0B",x"CD",x"C9", -- 0x2DD0
		x"6E",x"B7",x"06",x"09",x"28",x"0E",x"3D",x"18", -- 0x2DD8
		x"0A",x"CD",x"C9",x"6E",x"FE",x"09",x"06",x"00", -- 0x2DE0
		x"28",x"02",x"3C",x"47",x"78",x"81",x"32",x"96", -- 0x2DE8
		x"E9",x"CD",x"C9",x"6E",x"E6",x"0F",x"07",x"07", -- 0x2DF0
		x"07",x"07",x"C6",x"2C",x"6F",x"26",x"C4",x"78", -- 0x2DF8
		x"B7",x"28",x"07",x"7C",x"D6",x"10",x"67",x"05", -- 0x2E00
		x"18",x"F7",x"22",x"02",x"EB",x"3A",x"A4",x"E0", -- 0x2E08
		x"B7",x"CA",x"7A",x"6E",x"3D",x"32",x"A4",x"E0", -- 0x2E10
		x"C3",x"7A",x"6E",x"AF",x"32",x"A3",x"E0",x"32", -- 0x2E18
		x"A0",x"E0",x"21",x"A4",x"E0",x"7E",x"B7",x"28", -- 0x2E20
		x"04",x"35",x"C3",x"7A",x"6E",x"36",x"04",x"3A", -- 0x2E28
		x"96",x"E9",x"FE",x"25",x"38",x"24",x"20",x"04", -- 0x2E30
		x"3E",x"30",x"18",x"20",x"FE",x"26",x"20",x"59", -- 0x2E38
		x"3A",x"9B",x"E9",x"B7",x"28",x"34",x"3D",x"32", -- 0x2E40
		x"9B",x"E9",x"2A",x"90",x"E9",x"01",x"E0",x"FF", -- 0x2E48
		x"09",x"22",x"90",x"E9",x"36",x"30",x"DD",x"2B", -- 0x2E50
		x"18",x"20",x"C6",x"0A",x"2A",x"90",x"E9",x"77", -- 0x2E58
		x"DD",x"77",x"05",x"DD",x"23",x"01",x"20",x"00", -- 0x2E60
		x"09",x"22",x"90",x"E9",x"06",x"02",x"DF",x"3A", -- 0x2E68
		x"9B",x"E9",x"3C",x"32",x"9B",x"E9",x"FE",x"08", -- 0x2E70
		x"30",x"1F",x"06",x"02",x"DF",x"21",x"93",x"E9", -- 0x2E78
		x"35",x"C2",x"6C",x"6D",x"36",x"1E",x"11",x"95", -- 0x2E80
		x"E9",x"21",x"C4",x"78",x"06",x"02",x"CD",x"0E", -- 0x2E88
		x"02",x"2A",x"94",x"E9",x"7D",x"B4",x"C2",x"6C", -- 0x2E90
		x"6D",x"3E",x"03",x"32",x"9B",x"E9",x"DD",x"E5", -- 0x2E98
		x"E1",x"7D",x"E6",x"F8",x"C6",x"05",x"6F",x"06", -- 0x2EA0
		x"08",x"3E",x"30",x"BE",x"C0",x"23",x"10",x"FB", -- 0x2EA8
		x"2B",x"36",x"16",x"2B",x"36",x"18",x"2B",x"36", -- 0x2EB0
		x"0C",x"2B",x"36",x"19",x"2B",x"36",x"0A",x"2B", -- 0x2EB8
		x"36",x"0C",x"2B",x"36",x"30",x"2B",x"36",x"38", -- 0x2EC0
		x"C9",x"01",x"00",x"00",x"FE",x"0A",x"D8",x"D6", -- 0x2EC8
		x"0A",x"04",x"08",x"79",x"C6",x"0A",x"4F",x"08", -- 0x2ED0
		x"18",x"F2",x"06",x"9E",x"DF",x"3A",x"9B",x"E9", -- 0x2ED8
		x"FE",x"03",x"20",x"F6",x"3A",x"BF",x"EF",x"32", -- 0x2EE0
		x"A5",x"E9",x"F7",x"CD",x"0E",x"6F",x"CD",x"28", -- 0x2EE8
		x"6F",x"3A",x"92",x"E9",x"B7",x"20",x"01",x"2C", -- 0x2EF0
		x"11",x"C7",x"78",x"CD",x"48",x"6F",x"D9",x"21", -- 0x2EF8
		x"4E",x"D4",x"4F",x"06",x"1E",x"CD",x"49",x"02", -- 0x2F00
		x"D9",x"CD",x"34",x"6F",x"18",x"ED",x"3A",x"92", -- 0x2F08
		x"E9",x"4F",x"11",x"05",x"00",x"79",x"BB",x"38", -- 0x2F10
		x"07",x"93",x"4F",x"7A",x"83",x"57",x"18",x"F5", -- 0x2F18
		x"32",x"99",x"E9",x"7A",x"32",x"9A",x"E9",x"C9", -- 0x2F20
		x"3A",x"99",x"E9",x"07",x"4F",x"21",x"4A",x"D4", -- 0x2F28
		x"7D",x"91",x"6F",x"C9",x"C5",x"E5",x"CD",x"48", -- 0x2F30
		x"6F",x"D5",x"4F",x"06",x"1E",x"CD",x"49",x"02", -- 0x2F38
		x"D1",x"13",x"E1",x"06",x"04",x"DF",x"C1",x"C9", -- 0x2F40
		x"1A",x"FE",x"FF",x"C0",x"11",x"C7",x"78",x"1A", -- 0x2F48
		x"C9",x"3E",x"01",x"32",x"C7",x"E0",x"DD",x"21", -- 0x2F50
		x"A0",x"A2",x"CD",x"CC",x"2C",x"CD",x"88",x"25", -- 0x2F58
		x"CD",x"6C",x"24",x"21",x"5D",x"E1",x"11",x"6C", -- 0x2F60
		x"E7",x"01",x"03",x"00",x"ED",x"B0",x"CD",x"C1", -- 0x2F68
		x"24",x"3A",x"74",x"E7",x"21",x"78",x"E7",x"CD", -- 0x2F70
		x"BE",x"23",x"21",x"C0",x"E9",x"4E",x"3A",x"74", -- 0x2F78
		x"E7",x"B9",x"38",x"01",x"77",x"79",x"21",x"7B", -- 0x2F80
		x"E7",x"CD",x"BE",x"23",x"CD",x"ED",x"23",x"21", -- 0x2F88
		x"BF",x"A5",x"CD",x"70",x"23",x"21",x"77",x"D2", -- 0x2F90
		x"11",x"60",x"E7",x"06",x"08",x"CD",x"96",x"23", -- 0x2F98
		x"06",x"0A",x"DF",x"0E",x"1B",x"CD",x"78",x"11", -- 0x2FA0
		x"06",x"28",x"DF",x"21",x"F3",x"A5",x"CD",x"70", -- 0x2FA8
		x"23",x"21",x"F4",x"D2",x"11",x"78",x"E7",x"06", -- 0x2FB0
		x"03",x"CD",x"96",x"23",x"06",x"01",x"3E",x"29", -- 0x2FB8
		x"CD",x"B1",x"23",x"06",x"0A",x"DF",x"0E",x"1B", -- 0x2FC0
		x"CD",x"78",x"11",x"06",x"28",x"DF",x"21",x"E3", -- 0x2FC8
		x"A5",x"CD",x"70",x"23",x"21",x"F1",x"D2",x"11", -- 0x2FD0
		x"7B",x"E7",x"06",x"03",x"CD",x"96",x"23",x"06", -- 0x2FD8
		x"01",x"3E",x"29",x"CD",x"B1",x"23",x"06",x"0A", -- 0x2FE0
		x"DF",x"0E",x"1B",x"CD",x"78",x"11",x"06",x"28", -- 0x2FE8
		x"DF",x"21",x"A6",x"E9",x"CB",x"C6",x"F7",x"AF", -- 0x2FF0
		x"32",x"C7",x"EB",x"32",x"A6",x"E9",x"CD",x"E7", -- 0x2FF8
		x"2C",x"CD",x"A7",x"02",x"CD",x"D0",x"70",x"0E", -- 0x3000
		x"00",x"CD",x"78",x"11",x"0E",x"0B",x"CD",x"78", -- 0x3008
		x"11",x"0E",x"10",x"CD",x"78",x"11",x"0E",x"0F", -- 0x3010
		x"CD",x"78",x"11",x"DD",x"21",x"A0",x"A2",x"CD", -- 0x3018
		x"CC",x"2C",x"3E",x"05",x"01",x"51",x"6F",x"FF", -- 0x3020
		x"06",x"08",x"DF",x"3A",x"A6",x"E9",x"0F",x"30", -- 0x3028
		x"F7",x"06",x"28",x"DF",x"16",x"80",x"21",x"10", -- 0x3030
		x"D8",x"01",x"10",x"20",x"CD",x"53",x"02",x"16", -- 0x3038
		x"F8",x"21",x"00",x"D8",x"01",x"10",x"20",x"CD", -- 0x3040
		x"53",x"02",x"CD",x"D0",x"70",x"DD",x"21",x"7C", -- 0x3048
		x"A2",x"CD",x"CC",x"2C",x"3E",x"01",x"01",x"F2", -- 0x3050
		x"70",x"FF",x"21",x"85",x"A6",x"CD",x"70",x"23", -- 0x3058
		x"CD",x"E6",x"70",x"21",x"52",x"D1",x"06",x"0D", -- 0x3060
		x"11",x"12",x"A6",x"CD",x"96",x"23",x"CD",x"E6", -- 0x3068
		x"70",x"21",x"96",x"A6",x"CD",x"70",x"23",x"CD", -- 0x3070
		x"E6",x"70",x"21",x"CF",x"70",x"CD",x"D1",x"12", -- 0x3078
		x"21",x"8B",x"D1",x"11",x"49",x"A5",x"06",x"09", -- 0x3080
		x"CD",x"96",x"23",x"CD",x"E6",x"70",x"21",x"A9", -- 0x3088
		x"A6",x"CD",x"70",x"23",x"CD",x"E6",x"70",x"21", -- 0x3090
		x"C1",x"A6",x"CD",x"70",x"23",x"CD",x"E6",x"70", -- 0x3098
		x"21",x"C4",x"70",x"11",x"00",x"EB",x"01",x"04", -- 0x30A0
		x"00",x"ED",x"B0",x"06",x"00",x"DF",x"06",x"3C", -- 0x30A8
		x"DF",x"3E",x"01",x"EF",x"AF",x"32",x"01",x"E1", -- 0x30B0
		x"32",x"64",x"E1",x"32",x"1F",x"E1",x"32",x"07", -- 0x30B8
		x"EC",x"C3",x"96",x"69",x"D0",x"83",x"60",x"10", -- 0x30C0
		x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C8
		x"21",x"41",x"D0",x"01",x"1D",x"1C",x"16",x"30", -- 0x30D0
		x"CD",x"53",x"02",x"21",x"40",x"D4",x"01",x"1E", -- 0x30D8
		x"1C",x"16",x"00",x"C3",x"53",x"02",x"06",x"0A", -- 0x30E0
		x"DF",x"0E",x"1B",x"CD",x"78",x"11",x"06",x"28", -- 0x30E8
		x"DF",x"C9",x"21",x"50",x"D4",x"11",x"C7",x"78", -- 0x30F0
		x"CD",x"48",x"6F",x"CD",x"34",x"6F",x"18",x"F8", -- 0x30F8
		x"00",x"0D",x"22",x"D1",x"38",x"30",x"01",x"09", -- 0x3100
		x"08",x"04",x"30",x"0C",x"0A",x"19",x"0C",x"18", -- 0x3108
		x"16",x"00",x"ED",x"4B",x"64",x"EC",x"C5",x"DF", -- 0x3110
		x"C1",x"0D",x"20",x"FA",x"2A",x"60",x"EC",x"ED", -- 0x3118
		x"4B",x"62",x"EC",x"3A",x"BF",x"EF",x"0F",x"0F", -- 0x3120
		x"E6",x"FC",x"47",x"AE",x"23",x"0D",x"20",x"FB", -- 0x3128
		x"10",x"F9",x"47",x"3A",x"1C",x"00",x"B8",x"28", -- 0x3130
		x"2F",x"3A",x"BF",x"EF",x"47",x"C5",x"06",x"00", -- 0x3138
		x"DF",x"C1",x"10",x"F9",x"21",x"40",x"D0",x"01", -- 0x3140
		x"04",x"1C",x"16",x"30",x"CD",x"53",x"02",x"21", -- 0x3148
		x"40",x"D4",x"01",x"04",x"1C",x"16",x"16",x"CD", -- 0x3150
		x"53",x"02",x"21",x"00",x"71",x"CD",x"22",x"02", -- 0x3158
		x"21",x"69",x"71",x"CD",x"22",x"02",x"F3",x"76", -- 0x3160
		x"F7",x"00",x"19",x"83",x"D0",x"1B",x"18",x"16", -- 0x3168
		x"30",x"0E",x"1B",x"1B",x"18",x"1B",x"30",x"28", -- 0x3170
		x"30",x"0C",x"11",x"0E",x"0C",x"14",x"30",x"0A", -- 0x3178
		x"10",x"0A",x"12",x"17",x"30",x"28",x"00",x"00", -- 0x3180
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3188
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3190
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3198
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F8
		x"20",x"14",x"40",x"11",x"80",x"12",x"18",x"11", -- 0x3200
		x"04",x"12",x"04",x"02",x"04",x"12",x"04",x"02", -- 0x3208
		x"04",x"10",x"04",x"00",x"04",x"10",x"04",x"00", -- 0x3210
		x"04",x"10",x"04",x"00",x"04",x"10",x"04",x"00", -- 0x3218
		x"03",x"10",x"03",x"00",x"03",x"10",x"03",x"00", -- 0x3220
		x"03",x"12",x"03",x"02",x"03",x"12",x"03",x"02", -- 0x3228
		x"03",x"01",x"03",x"11",x"03",x"01",x"03",x"11", -- 0x3230
		x"03",x"00",x"03",x"10",x"03",x"00",x"03",x"10", -- 0x3238
		x"03",x"00",x"03",x"10",x"03",x"00",x"03",x"10", -- 0x3240
		x"03",x"08",x"20",x"18",x"08",x"10",x"10",x"11", -- 0x3248
		x"10",x"12",x"04",x"04",x"04",x"14",x"04",x"04", -- 0x3250
		x"04",x"14",x"04",x"04",x"04",x"14",x"04",x"04", -- 0x3258
		x"04",x"14",x"04",x"04",x"04",x"14",x"04",x"04", -- 0x3260
		x"30",x"18",x"04",x"04",x"04",x"14",x"04",x"04", -- 0x3268
		x"04",x"14",x"04",x"04",x"04",x"14",x"04",x"04", -- 0x3270
		x"04",x"14",x"04",x"04",x"04",x"14",x"04",x"04", -- 0x3278
		x"38",x"18",x"04",x"00",x"40",x"31",x"40",x"12", -- 0x3280
		x"20",x"14",x"10",x"19",x"04",x"00",x"04",x"11", -- 0x3288
		x"04",x"00",x"04",x"11",x"04",x"00",x"04",x"11", -- 0x3290
		x"04",x"00",x"04",x"11",x"04",x"00",x"04",x"11", -- 0x3298
		x"04",x"00",x"04",x"11",x"04",x"00",x"04",x"11", -- 0x32A0
		x"04",x"12",x"06",x"02",x"06",x"12",x"06",x"02", -- 0x32A8
		x"06",x"12",x"06",x"00",x"06",x"10",x"06",x"00", -- 0x32B0
		x"06",x"10",x"06",x"00",x"06",x"10",x"06",x"00", -- 0x32B8
		x"30",x"10",x"08",x"10",x"08",x"00",x"08",x"10", -- 0x32C0
		x"08",x"00",x"08",x"10",x"08",x"00",x"08",x"10", -- 0x32C8
		x"08",x"00",x"08",x"10",x"20",x"15",x"08",x"12", -- 0x32D0
		x"05",x"02",x"03",x"02",x"03",x"00",x"03",x"02", -- 0x32D8
		x"03",x"00",x"04",x"10",x"04",x"00",x"04",x"10", -- 0x32E0
		x"04",x"00",x"04",x"10",x"04",x"00",x"04",x"10", -- 0x32E8
		x"04",x"00",x"04",x"10",x"04",x"00",x"04",x"10", -- 0x32F0
		x"04",x"00",x"04",x"10",x"04",x"00",x"30",x"14", -- 0x32F8
		x"80",x"10",x"40",x"19",x"30",x"12",x"20",x"10", -- 0x3300
		x"10",x"08",x"01",x"08",x"11",x"08",x"01",x"08", -- 0x3308
		x"04",x"11",x"04",x"01",x"04",x"11",x"20",x"01", -- 0x3310
		x"80",x"14",x"20",x"14",x"40",x"11",x"60",x"1A", -- 0x3318
		x"04",x"10",x"04",x"00",x"04",x"10",x"04",x"00", -- 0x3320
		x"04",x"10",x"04",x"00",x"04",x"10",x"04",x"00", -- 0x3328
		x"20",x"15",x"20",x"11",x"08",x"10",x"08",x"00", -- 0x3330
		x"08",x"10",x"08",x"00",x"08",x"10",x"08",x"00", -- 0x3338
		x"50",x"16",x"20",x"1A",x"60",x"11",x"10",x"12", -- 0x3340
		x"30",x"10",x"20",x"14",x"30",x"11",x"18",x"1A", -- 0x3348
		x"30",x"18",x"40",x"16",x"30",x"15",x"30",x"18", -- 0x3350
		x"50",x"16",x"40",x"18",x"00",x"FF",x"10",x"10", -- 0x3358
		x"11",x"40",x"12",x"10",x"18",x"30",x"15",x"48", -- 0x3360
		x"19",x"10",x"04",x"03",x"12",x"03",x"02",x"03", -- 0x3368
		x"12",x"03",x"02",x"03",x"12",x"03",x"02",x"05", -- 0x3370
		x"10",x"05",x"00",x"05",x"10",x"05",x"00",x"05", -- 0x3378
		x"10",x"05",x"00",x"05",x"10",x"05",x"00",x"05", -- 0x3380
		x"10",x"05",x"00",x"05",x"10",x"05",x"00",x"05", -- 0x3388
		x"10",x"05",x"00",x"05",x"10",x"05",x"00",x"05", -- 0x3390
		x"10",x"05",x"00",x"05",x"10",x"70",x"00",x"40", -- 0x3398
		x"18",x"60",x"14",x"03",x"10",x"30",x"12",x"60", -- 0x33A0
		x"11",x"18",x"18",x"20",x"1A",x"30",x"16",x"10", -- 0x33A8
		x"15",x"10",x"18",x"18",x"19",x"03",x"08",x"03", -- 0x33B0
		x"10",x"03",x"00",x"03",x"10",x"03",x"08",x"03", -- 0x33B8
		x"10",x"03",x"00",x"03",x"10",x"03",x"08",x"03", -- 0x33C0
		x"10",x"03",x"00",x"03",x"10",x"03",x"00",x"03", -- 0x33C8
		x"11",x"03",x"00",x"03",x"11",x"03",x"00",x"03", -- 0x33D0
		x"11",x"03",x"00",x"03",x"1A",x"03",x"00",x"03", -- 0x33D8
		x"1A",x"03",x"00",x"03",x"12",x"03",x"00",x"03", -- 0x33E0
		x"1A",x"03",x"00",x"03",x"12",x"03",x"00",x"03", -- 0x33E8
		x"12",x"03",x"00",x"03",x"12",x"03",x"00",x"03", -- 0x33F0
		x"10",x"03",x"01",x"03",x"10",x"03",x"02",x"03", -- 0x33F8
		x"1A",x"03",x"02",x"03",x"1A",x"03",x"00",x"03", -- 0x3400
		x"1A",x"03",x"00",x"03",x"1A",x"06",x"02",x"06", -- 0x3408
		x"10",x"06",x"00",x"06",x"10",x"06",x"00",x"06", -- 0x3410
		x"12",x"06",x"02",x"06",x"12",x"06",x"02",x"06", -- 0x3418
		x"12",x"06",x"02",x"06",x"12",x"30",x"15",x"06", -- 0x3420
		x"12",x"06",x"02",x"06",x"12",x"00",x"00",x"00", -- 0x3428
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3430
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3438
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3440
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3448
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3450
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3458
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3460
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3468
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3470
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3478
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3480
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3488
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3490
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3498
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3500
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3508
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3510
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3518
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3520
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3528
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3530
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3538
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3540
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3548
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3550
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3558
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3560
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3568
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3570
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3578
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3580
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3588
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3590
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3598
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3600
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3608
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3610
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3618
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3620
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3628
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3630
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3638
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3640
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3648
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3650
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3658
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3660
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3668
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3670
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3678
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3680
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3688
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3690
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3698
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3700
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3708
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3710
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3718
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3720
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3728
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3730
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3738
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3740
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3748
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3750
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3760
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3768
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3770
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3778
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3798
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F8
		x"6A",x"01",x"6A",x"01",x"6A",x"01",x"6A",x"01", -- 0x3800
		x"6A",x"01",x"6A",x"01",x"6A",x"01",x"6A",x"01", -- 0x3808
		x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"02", -- 0x3810
		x"00",x"02",x"00",x"00",x"00",x"02",x"00",x"00", -- 0x3818
		x"C4",x"00",x"D9",x"01",x"D9",x"01",x"C4",x"00", -- 0x3820
		x"C4",x"00",x"D9",x"01",x"D9",x"01",x"C4",x"00", -- 0x3828
		x"C4",x"00",x"D9",x"01",x"D9",x"01",x"C4",x"00", -- 0x3830
		x"C4",x"00",x"D9",x"01",x"D9",x"01",x"C4",x"00", -- 0x3838
		x"C5",x"01",x"C5",x"01",x"C5",x"01",x"C5",x"01", -- 0x3840
		x"C5",x"01",x"C5",x"01",x"C5",x"01",x"C5",x"01", -- 0x3848
		x"00",x"00",x"80",x"02",x"00",x"00",x"80",x"02", -- 0x3850
		x"80",x"02",x"00",x"00",x"80",x"02",x"00",x"00", -- 0x3858
		x"F5",x"00",x"4F",x"02",x"4F",x"02",x"F5",x"00", -- 0x3860
		x"F5",x"00",x"4F",x"02",x"4F",x"02",x"F5",x"00", -- 0x3868
		x"F5",x"00",x"4F",x"02",x"4F",x"02",x"F5",x"00", -- 0x3870
		x"F5",x"00",x"4F",x"02",x"4F",x"02",x"F5",x"00", -- 0x3878
		x"05",x"02",x"01",x"03",x"E8",x"E0",x"06",x"EA", -- 0x3880
		x"E2",x"08",x"EC",x"E4",x"08",x"EE",x"E6",x"08", -- 0x3888
		x"FC",x"F4",x"08",x"EE",x"E6",x"06",x"FC",x"F4", -- 0x3890
		x"08",x"FE",x"F6",x"08",x"00",x"00",x"00",x"04", -- 0x3898
		x"01",x"03",x"01",x"02",x"03",x"02",x"01",x"01", -- 0x38A0
		x"04",x"01",x"02",x"01",x"01",x"00",x"00",x"04", -- 0x38A8
		x"01",x"03",x"01",x"02",x"03",x"02",x"01",x"01", -- 0x38B0
		x"04",x"01",x"02",x"01",x"01",x"00",x"00",x"00", -- 0x38B8
		x"00",x"00",x"00",x"00",x"01",x"00",x"02",x"16", -- 0x38C0
		x"17",x"19",x"1A",x"1B",x"1C",x"1D",x"1E",x"12", -- 0x38C8
		x"11",x"14",x"15",x"FF",x"00",x"40",x"41",x"42", -- 0x38D0
		x"10",x"44",x"45",x"46",x"20",x"48",x"49",x"4A", -- 0x38D8
		x"30",x"4C",x"4D",x"4E",x"00",x"01",x"02",x"03", -- 0x38E0
		x"04",x"05",x"06",x"07",x"10",x"11",x"12",x"13", -- 0x38E8
		x"14",x"15",x"16",x"17",x"20",x"21",x"22",x"23", -- 0x38F0
		x"0B",x"25",x"26",x"27",x"30",x"31",x"32",x"33", -- 0x38F8
		x"1B",x"35",x"36",x"37",x"00",x"08",x"09",x"0A", -- 0x3900
		x"0B",x"0C",x"0D",x"0E",x"10",x"18",x"19",x"1A", -- 0x3908
		x"1B",x"1C",x"1D",x"1E",x"20",x"28",x"29",x"2A", -- 0x3910
		x"04",x"2C",x"2D",x"2E",x"30",x"38",x"39",x"3A", -- 0x3918
		x"14",x"3C",x"3D",x"3E",x"58",x"59",x"5A",x"5B", -- 0x3920
		x"5C",x"5D",x"5E",x"5F",x"50",x"51",x"52",x"53", -- 0x3928
		x"54",x"55",x"56",x"57",x"FF",x"FF",x"FF",x"FF", -- 0x3930
		x"FF",x"FF",x"FF",x"FF",x"58",x"78",x"79",x"7A", -- 0x3938
		x"7B",x"7C",x"7D",x"7E",x"FF",x"FF",x"FF",x"FF", -- 0x3940
		x"FF",x"FF",x"FF",x"FF",x"50",x"70",x"71",x"72", -- 0x3948
		x"73",x"74",x"75",x"76",x"68",x"69",x"6A",x"6B", -- 0x3950
		x"6C",x"6D",x"6E",x"6F",x"60",x"61",x"62",x"63", -- 0x3958
		x"64",x"65",x"66",x"67",x"68",x"70",x"71",x"72", -- 0x3960
		x"73",x"74",x"75",x"76",x"FF",x"FF",x"FF",x"FF", -- 0x3968
		x"FF",x"FF",x"FF",x"FF",x"60",x"78",x"79",x"7A", -- 0x3970
		x"7B",x"7C",x"7D",x"7E",x"FF",x"01",x"FF",x"FF", -- 0x3978
		x"01",x"01",x"01",x"FF",x"00",x"01",x"00",x"FF", -- 0x3980
		x"FF",x"00",x"01",x"00",x"94",x"79",x"98",x"79", -- 0x3988
		x"98",x"79",x"94",x"79",x"01",x"01",x"01",x"FF", -- 0x3990
		x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"A5", -- 0x3998
		x"79",x"4E",x"7A",x"1B",x"7B",x"01",x"40",x"FE", -- 0x39A0
		x"00",x"01",x"40",x"FF",x"00",x"01",x"40",x"FE", -- 0x39A8
		x"00",x"01",x"40",x"FF",x"00",x"01",x"40",x"FE", -- 0x39B0
		x"00",x"08",x"40",x"FF",x"00",x"02",x"41",x"FF", -- 0x39B8
		x"00",x"01",x"41",x"FF",x"01",x"01",x"41",x"FF", -- 0x39C0
		x"00",x"01",x"41",x"00",x"00",x"02",x"41",x"FF", -- 0x39C8
		x"00",x"01",x"41",x"FF",x"01",x"01",x"41",x"FF", -- 0x39D0
		x"00",x"01",x"41",x"00",x"00",x"02",x"41",x"FF", -- 0x39D8
		x"00",x"01",x"41",x"FF",x"01",x"01",x"41",x"FF", -- 0x39E0
		x"00",x"01",x"41",x"00",x"00",x"01",x"42",x"FF", -- 0x39E8
		x"01",x"01",x"42",x"00",x"00",x"01",x"42",x"FF", -- 0x39F0
		x"01",x"01",x"42",x"00",x"00",x"01",x"42",x"FF", -- 0x39F8
		x"01",x"01",x"42",x"00",x"00",x"01",x"42",x"FF", -- 0x3A00
		x"01",x"01",x"42",x"00",x"00",x"01",x"42",x"00", -- 0x3A08
		x"01",x"01",x"42",x"00",x"00",x"01",x"42",x"00", -- 0x3A10
		x"01",x"01",x"42",x"00",x"00",x"01",x"43",x"00", -- 0x3A18
		x"01",x"01",x"43",x"00",x"00",x"01",x"43",x"00", -- 0x3A20
		x"01",x"01",x"43",x"00",x"00",x"04",x"43",x"01", -- 0x3A28
		x"01",x"01",x"44",x"02",x"00",x"01",x"44",x"02", -- 0x3A30
		x"01",x"01",x"44",x"02",x"00",x"01",x"44",x"02", -- 0x3A38
		x"01",x"01",x"44",x"02",x"00",x"01",x"44",x"02", -- 0x3A40
		x"01",x"08",x"44",x"02",x"00",x"00",x"01",x"40", -- 0x3A48
		x"FE",x"01",x"01",x"40",x"FE",x"00",x"01",x"40", -- 0x3A50
		x"FE",x"01",x"01",x"40",x"FE",x"00",x"01",x"40", -- 0x3A58
		x"FE",x"01",x"01",x"40",x"FE",x"00",x"02",x"40", -- 0x3A60
		x"FE",x"01",x"01",x"41",x"FE",x"01",x"01",x"41", -- 0x3A68
		x"00",x"00",x"01",x"41",x"FE",x"01",x"01",x"41", -- 0x3A70
		x"00",x"00",x"01",x"41",x"FE",x"01",x"01",x"41", -- 0x3A78
		x"00",x"00",x"02",x"41",x"FF",x"01",x"01",x"41", -- 0x3A80
		x"FF",x"00",x"01",x"41",x"FF",x"01",x"01",x"41", -- 0x3A88
		x"FF",x"00",x"04",x"42",x"FF",x"01",x"01",x"42", -- 0x3A90
		x"00",x"01",x"01",x"42",x"FF",x"01",x"01",x"42", -- 0x3A98
		x"00",x"01",x"01",x"42",x"00",x"00",x"01",x"42", -- 0x3AA0
		x"00",x"01",x"01",x"42",x"00",x"00",x"01",x"42", -- 0x3AA8
		x"00",x"01",x"01",x"42",x"00",x"00",x"01",x"43", -- 0x3AB0
		x"00",x"01",x"01",x"43",x"00",x"00",x"01",x"43", -- 0x3AB8
		x"00",x"01",x"01",x"43",x"00",x"00",x"01",x"43", -- 0x3AC0
		x"01",x"01",x"01",x"43",x"00",x"01",x"04",x"44", -- 0x3AC8
		x"01",x"01",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3AD0
		x"00",x"00",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3AD8
		x"00",x"00",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3AE0
		x"00",x"00",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3AE8
		x"00",x"00",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3AF0
		x"00",x"00",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3AF8
		x"02",x"00",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3B00
		x"02",x"00",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3B08
		x"02",x"00",x"01",x"44",x"02",x"01",x"01",x"44", -- 0x3B10
		x"02",x"00",x"00",x"04",x"40",x"FE",x"01",x"01", -- 0x3B18
		x"40",x"FE",x"01",x"01",x"40",x"00",x"00",x"01", -- 0x3B20
		x"40",x"FE",x"01",x"01",x"40",x"00",x"00",x"01", -- 0x3B28
		x"40",x"FE",x"01",x"01",x"40",x"00",x"00",x"01", -- 0x3B30
		x"40",x"FE",x"01",x"01",x"40",x"00",x"00",x"03", -- 0x3B38
		x"41",x"FF",x"01",x"01",x"41",x"FF",x"00",x"03", -- 0x3B40
		x"41",x"FF",x"01",x"01",x"41",x"00",x"01",x"03", -- 0x3B48
		x"41",x"FF",x"01",x"01",x"42",x"FF",x"01",x"01", -- 0x3B50
		x"42",x"00",x"01",x"02",x"42",x"FF",x"01",x"01", -- 0x3B58
		x"42",x"00",x"01",x"01",x"42",x"FF",x"01",x"02", -- 0x3B60
		x"42",x"00",x"01",x"01",x"42",x"FF",x"01",x"03", -- 0x3B68
		x"42",x"00",x"01",x"03",x"43",x"00",x"01",x"01", -- 0x3B70
		x"43",x"01",x"01",x"02",x"43",x"00",x"01",x"01", -- 0x3B78
		x"43",x"01",x"01",x"01",x"43",x"00",x"01",x"01", -- 0x3B80
		x"43",x"01",x"01",x"01",x"43",x"00",x"01",x"01", -- 0x3B88
		x"43",x"01",x"01",x"03",x"44",x"01",x"01",x"01", -- 0x3B90
		x"44",x"00",x"01",x"03",x"44",x"01",x"01",x"01", -- 0x3B98
		x"44",x"01",x"00",x"03",x"44",x"01",x"01",x"01", -- 0x3BA0
		x"44",x"00",x"00",x"01",x"44",x"02",x"01",x"01", -- 0x3BA8
		x"44",x"00",x"00",x"01",x"44",x"02",x"01",x"01", -- 0x3BB0
		x"44",x"00",x"00",x"01",x"44",x"02",x"01",x"01", -- 0x3BB8
		x"44",x"00",x"00",x"01",x"44",x"02",x"01",x"04", -- 0x3BC0
		x"44",x"02",x"01",x"00",x"01",x"FE",x"01",x"01", -- 0x3BC8
		x"FE",x"00",x"01",x"FE",x"01",x"01",x"FE",x"00", -- 0x3BD0
		x"01",x"FE",x"01",x"01",x"FE",x"00",x"01",x"FE", -- 0x3BD8
		x"01",x"01",x"FE",x"00",x"03",x"FE",x"01",x"01", -- 0x3BE0
		x"FE",x"00",x"03",x"FE",x"01",x"01",x"FE",x"02", -- 0x3BE8
		x"03",x"FE",x"01",x"11",x"FE",x"02",x"01",x"FF", -- 0x3BF0
		x"02",x"02",x"FE",x"02",x"01",x"FF",x"02",x"01", -- 0x3BF8
		x"FE",x"02",x"01",x"FF",x"02",x"01",x"FE",x"02", -- 0x3C00
		x"01",x"FF",x"02",x"01",x"FE",x"02",x"01",x"FF", -- 0x3C08
		x"02",x"01",x"FE",x"02",x"01",x"FF",x"02",x"01", -- 0x3C10
		x"FE",x"02",x"01",x"FF",x"02",x"01",x"FE",x"02", -- 0x3C18
		x"63",x"FF",x"02",x"00",x"00",x"02",x"00",x"FE", -- 0x3C20
		x"FE",x"00",x"02",x"00",x"FE",x"01",x"FE",x"FF", -- 0x3C28
		x"FF",x"FE",x"01",x"FE",x"00",x"01",x"FF",x"02", -- 0x3C30
		x"03",x"04",x"FF",x"05",x"06",x"07",x"00",x"02", -- 0x3C38
		x"03",x"01",x"03",x"00",x"01",x"02",x"00",x"40", -- 0x3C40
		x"41",x"42",x"10",x"44",x"45",x"46",x"20",x"48", -- 0x3C48
		x"49",x"4A",x"30",x"4C",x"4D",x"4E",x"76",x"7C", -- 0x3C50
		x"8E",x"7C",x"92",x"7C",x"96",x"7C",x"7C",x"7C", -- 0x3C58
		x"9A",x"7C",x"9E",x"7C",x"A2",x"7C",x"82",x"7C", -- 0x3C60
		x"A6",x"7C",x"AA",x"7C",x"AE",x"7C",x"88",x"7C", -- 0x3C68
		x"B2",x"7C",x"B6",x"7C",x"BA",x"7C",x"07",x"02", -- 0x3C70
		x"03",x"0D",x"0F",x"FF",x"05",x"01",x"03",x"0A", -- 0x3C78
		x"0E",x"FF",x"06",x"00",x"01",x"09",x"0B",x"FF", -- 0x3C80
		x"04",x"02",x"00",x"08",x"0C",x"FF",x"07",x"0F", -- 0x3C88
		x"03",x"FF",x"03",x"0E",x"0F",x"FF",x"03",x"0E", -- 0x3C90
		x"05",x"FF",x"05",x"0A",x"01",x"FF",x"01",x"0A", -- 0x3C98
		x"0B",x"FF",x"01",x"0B",x"06",x"FF",x"06",x"09", -- 0x3CA0
		x"00",x"FF",x"00",x"08",x"09",x"FF",x"00",x"08", -- 0x3CA8
		x"04",x"FF",x"04",x"0C",x"02",x"FF",x"02",x"0C", -- 0x3CB0
		x"0D",x"FF",x"02",x"0D",x"07",x"FF",x"0C",x"00", -- 0x3CB8
		x"0B",x"FD",x"0B",x"FB",x"09",x"FB",x"06",x"FA", -- 0x3CC0
		x"03",x"FB",x"01",x"FB",x"01",x"FD",x"00",x"00", -- 0x3CC8
		x"01",x"03",x"01",x"05",x"03",x"05",x"06",x"06", -- 0x3CD0
		x"09",x"05",x"0B",x"05",x"0B",x"03",x"17",x"07", -- 0x3CD8
		x"17",x"03",x"15",x"02",x"13",x"00",x"0F",x"00", -- 0x3CE0
		x"0C",x"00",x"09",x"01",x"08",x"04",x"08",x"07", -- 0x3CE8
		x"08",x"0C",x"0A",x"0E",x"0D",x"0F",x"0F",x"0F", -- 0x3CF0
		x"13",x"10",x"15",x"0D",x"17",x"0A",x"17",x"07", -- 0x3CF8
		x"17",x"03",x"15",x"02",x"13",x"00",x"0F",x"00", -- 0x3D00
		x"0C",x"00",x"09",x"01",x"08",x"04",x"18",x"60", -- 0x3D08
		x"10",x"60",x"04",x"A0",x"00",x"20",x"1A",x"60", -- 0x3D10
		x"12",x"60",x"08",x"A0",x"01",x"20",x"1E",x"60", -- 0x3D18
		x"1C",x"60",x"0C",x"A0",x"01",x"20",x"F0",x"00", -- 0x3D20
		x"22",x"60",x"14",x"A0",x"02",x"20",x"F0",x"00", -- 0x3D28
		x"28",x"60",x"24",x"A0",x"F0",x"00",x"F0",x"00", -- 0x3D30
		x"2A",x"60",x"2C",x"A0",x"F0",x"00",x"F0",x"00", -- 0x3D38
		x"32",x"60",x"34",x"A0",x"F0",x"00",x"18",x"60", -- 0x3D40
		x"58",x"60",x"40",x"A0",x"00",x"20",x"18",x"60", -- 0x3D48
		x"5A",x"60",x"44",x"A0",x"00",x"20",x"18",x"60", -- 0x3D50
		x"5C",x"60",x"48",x"A0",x"00",x"20",x"18",x"60", -- 0x3D58
		x"5E",x"60",x"4C",x"A0",x"00",x"20",x"18",x"60", -- 0x3D60
		x"60",x"60",x"50",x"A0",x"00",x"20",x"18",x"60", -- 0x3D68
		x"62",x"60",x"54",x"A0",x"00",x"20",x"31",x"08", -- 0x3D70
		x"15",x"06",x"15",x"09",x"06",x"08",x"8E",x"7D", -- 0x3D78
		x"96",x"7D",x"9E",x"7D",x"A6",x"7D",x"AE",x"7D", -- 0x3D80
		x"B6",x"7D",x"BE",x"7D",x"C6",x"7D",x"00",x"04", -- 0x3D88
		x"07",x"00",x"04",x"07",x"00",x"04",x"01",x"05", -- 0x3D90
		x"06",x"01",x"05",x"06",x"01",x"05",x"02",x"04", -- 0x3D98
		x"06",x"02",x"04",x"06",x"02",x"04",x"03",x"05", -- 0x3DA0
		x"07",x"03",x"05",x"07",x"03",x"05",x"04",x"02", -- 0x3DA8
		x"00",x"04",x"02",x"00",x"04",x"02",x"05",x"01", -- 0x3DB0
		x"03",x"05",x"01",x"03",x"05",x"01",x"06",x"01", -- 0x3DB8
		x"02",x"06",x"01",x"02",x"06",x"01",x"07",x"00", -- 0x3DC0
		x"03",x"07",x"00",x"03",x"07",x"00",x"10",x"00", -- 0x3DC8
		x"10",x"30",x"08",x"40",x"10",x"50",x"10",x"60", -- 0x3DD0
		x"06",x"80",x"00",x"10",x"80",x"10",x"70",x"08", -- 0x3DD8
		x"60",x"10",x"40",x"10",x"20",x"06",x"00",x"00", -- 0x3DE0
		x"08",x"80",x"0A",x"00",x"08",x"40",x"0A",x"30", -- 0x3DE8
		x"08",x"00",x"00",x"08",x"00",x"0A",x"30",x"08", -- 0x3DF0
		x"50",x"0A",x"60",x"02",x"70",x"06",x"80",x"00", -- 0x3DF8
		x"18",x"7E",x"27",x"7E",x"3A",x"7E",x"49",x"7E", -- 0x3E00
		x"66",x"7E",x"7B",x"7E",x"57",x"7E",x"18",x"7E", -- 0x3E08
		x"70",x"7E",x"27",x"7E",x"83",x"7E",x"3A",x"7E", -- 0x3E10
		x"08",x"30",x"08",x"60",x"08",x"70",x"60",x"80", -- 0x3E18
		x"08",x"70",x"08",x"60",x"08",x"30",x"00",x"08", -- 0x3E20
		x"20",x"08",x"60",x"08",x"60",x"08",x"70",x"18", -- 0x3E28
		x"80",x"08",x"70",x"08",x"60",x"08",x"60",x"08", -- 0x3E30
		x"20",x"00",x"08",x"10",x"08",x"20",x"08",x"60", -- 0x3E38
		x"0C",x"70",x"08",x"60",x"08",x"20",x"08",x"10", -- 0x3E40
		x"00",x"08",x"00",x"18",x"10",x"08",x"20",x"08", -- 0x3E48
		x"30",x"08",x"40",x"08",x"50",x"08",x"70",x"08", -- 0x3E50
		x"70",x"08",x"50",x"08",x"40",x"08",x"30",x"08", -- 0x3E58
		x"20",x"18",x"10",x"08",x"00",x"00",x"0C",x"18", -- 0x3E60
		x"08",x"40",x"08",x"40",x"08",x"70",x"08",x"80", -- 0x3E68
		x"08",x"80",x"08",x"70",x"08",x"40",x"08",x"40", -- 0x3E70
		x"0C",x"18",x"00",x"06",x"28",x"08",x"60",x"08", -- 0x3E78
		x"80",x"08",x"80",x"08",x"80",x"08",x"80",x"08", -- 0x3E80
		x"60",x"06",x"28",x"00",x"47",x"B1",x"02",x"00", -- 0x3E88
		x"47",x"D7",x"02",x"05",x"4B",x"B1",x"03",x"00", -- 0x3E90
		x"4B",x"D7",x"03",x"05",x"4F",x"B1",x"04",x"00", -- 0x3E98
		x"4F",x"D7",x"04",x"05",x"B2",x"B1",x"05",x"00", -- 0x3EA0
		x"B2",x"D7",x"05",x"05",x"7F",x"B1",x"06",x"00", -- 0x3EA8
		x"7F",x"D7",x"06",x"05",x"8E",x"B1",x"07",x"00", -- 0x3EB0
		x"8E",x"D7",x"07",x"05",x"8F",x"B1",x"08",x"00", -- 0x3EB8
		x"8F",x"D7",x"08",x"05",x"77",x"B1",x"09",x"00", -- 0x3EC0
		x"00",x"00",x"F0",x"10",x"00",x"20",x"F0",x"30", -- 0x3EC8
		x"B0",x"40",x"D0",x"40",x"D0",x"50",x"00",x"60", -- 0x3ED0
		x"10",x"00",x"10",x"10",x"10",x"20",x"10",x"30", -- 0x3ED8
		x"10",x"40",x"50",x"40",x"10",x"50",x"10",x"60", -- 0x3EE0
		x"C0",x"2E",x"C2",x"6E",x"C1",x"2E",x"C6",x"6E", -- 0x3EE8
		x"CC",x"6E",x"C8",x"AE",x"D0",x"AE",x"CE",x"2E", -- 0x3EF0
		x"D6",x"2E",x"D4",x"6E",x"D7",x"2E",x"D8",x"6E", -- 0x3EF8
		x"DC",x"AE",x"E4",x"6E",x"E0",x"AE",x"CF",x"2E", -- 0x3F00
		x"40",x"20",x"20",x"30",x"10",x"40",x"50",x"40", -- 0x3F08
		x"00",x"10",x"21",x"80",x"41",x"00",x"A0",x"20", -- 0x3F10
		x"20",x"10",x"04",x"00",x"10",x"21",x"00",x"50", -- 0x3F18
		x"41",x"10",x"21",x"04",x"00",x"20",x"10",x"00", -- 0x3F20
		x"66",x"08",x"28",x"02",x"28",x"0C",x"0E",x"08", -- 0x3F28
		x"3D",x"08",x"40",x"E2",x"40",x"28",x"02",x"07", -- 0x3F30
		x"01",x"01",x"01",x"05",x"01",x"03",x"02",x"06", -- 0x3F38
		x"00",x"00",x"00",x"04",x"00",x"03",x"00",x"01", -- 0x3F40
		x"00",x"FF",x"FF",x"00",x"01",x"00",x"01",x"01", -- 0x3F48
		x"01",x"FF",x"FF",x"01",x"FF",x"FF",x"04",x"08", -- 0x3F50
		x"40",x"08",x"48",x"E8",x"48",x"28",x"20",x"08", -- 0x3F58
		x"05",x"06",x"58",x"08",x"10",x"08",x"30",x"00", -- 0x3F60
		x"44",x"40",x"48",x"D8",x"06",x"05",x"4C",x"F8", -- 0x3F68
		x"4C",x"E8",x"4C",x"D8",x"4C",x"18",x"4C",x"28", -- 0x3F70
		x"4C",x"38",x"04",x"03",x"38",x"08",x"44",x"D0", -- 0x3F78
		x"54",x"10",x"14",x"14",x"04",x"03",x"18",x"80", -- 0x3F80
		x"3C",x"24",x"40",x"E8",x"48",x"20",x"04",x"03", -- 0x3F88
		x"28",x"08",x"44",x"C0",x"30",x"10",x"44",x"38", -- 0x3F90
		x"04",x"03",x"4C",x"00",x"3C",x"28",x"10",x"08", -- 0x3F98
		x"58",x"10",x"04",x"03",x"38",x"F8",x"48",x"48", -- 0x3FA0
		x"48",x"E8",x"40",x"08",x"04",x"07",x"18",x"10", -- 0x3FA8
		x"50",x"F0",x"38",x"28",x"48",x"C8",x"0C",x"03", -- 0x3FB0
		x"10",x"08",x"18",x"04",x"14",x"14",x"28",x"08", -- 0x3FB8
		x"44",x"D0",x"4C",x"E0",x"40",x"F8",x"50",x"08", -- 0x3FC0
		x"4C",x"18",x"44",x"30",x"4C",x"48",x"60",x"08", -- 0x3FC8
		x"00",x"DB",x"7F",x"E5",x"7F",x"EF",x"7F",x"F9", -- 0x3FD0
		x"7F",x"03",x"80",x"0D",x"80",x"0D",x"80",x"0D", -- 0x3FD8
		x"80",x"0D",x"80",x"0D",x"80",x"12",x"81",x"12", -- 0x3FE0
		x"81",x"12",x"81",x"12",x"81",x"12",x"81",x"9F", -- 0x3FE8
		x"82",x"9F",x"82",x"9F",x"82",x"9F",x"82",x"9F", -- 0x3FF0
		x"82",x"E4",x"82",x"25",x"83",x"AA",x"83",x"2F"  -- 0x3FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
