-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_A4 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_A4 is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"DC",x"B6",x"AF",x"8E",x"88",x"56",x"8D",x"C6", -- 0x0000
		x"84",x"81",x"53",x"A2",x"91",x"C5",x"CE",x"DE", -- 0x0008
		x"CB",x"D1",x"7A",x"BF",x"7E",x"FB",x"7B",x"F5", -- 0x0010
		x"72",x"2E",x"0D",x"20",x"91",x"06",x"A9",x"CF", -- 0x0018
		x"55",x"AB",x"AA",x"55",x"55",x"AA",x"52",x"D5", -- 0x0020
		x"FB",x"FD",x"BE",x"3E",x"BE",x"17",x"87",x"5F", -- 0x0028
		x"4B",x"51",x"B2",x"AA",x"5C",x"55",x"BB",x"AA", -- 0x0030
		x"65",x"75",x"DA",x"AA",x"99",x"54",x"54",x"AA", -- 0x0038
		x"EF",x"4F",x"9B",x"D5",x"B0",x"49",x"03",x"8F", -- 0x0040
		x"EA",x"55",x"DD",x"3A",x"09",x"91",x"C2",x"6E", -- 0x0048
		x"CB",x"D5",x"56",x"0B",x"DC",x"F7",x"FB",x"FA", -- 0x0050
		x"F5",x"FD",x"FE",x"7E",x"45",x"8E",x"18",x"F8", -- 0x0058
		x"FF",x"DF",x"0D",x"54",x"89",x"60",x"7E",x"1F", -- 0x0060
		x"2A",x"84",x"42",x"A5",x"F3",x"ED",x"DE",x"E6", -- 0x0068
		x"53",x"11",x"B2",x"6A",x"FC",x"F5",x"7B",x"9A", -- 0x0070
		x"25",x"35",x"5A",x"EB",x"FA",x"F6",x"F6",x"FA", -- 0x0078
		x"B3",x"46",x"05",x"10",x"D8",x"7D",x"67",x"2F", -- 0x0080
		x"85",x"C0",x"05",x"6B",x"42",x"05",x"0D",x"0C", -- 0x0088
		x"F8",x"DD",x"BA",x"6B",x"EC",x"D7",x"3B",x"AA", -- 0x0090
		x"C5",x"FD",x"DE",x"AA",x"99",x"54",x"54",x"AA", -- 0x0098
		x"19",x"13",x"FA",x"FD",x"BD",x"6A",x"96",x"15", -- 0x00A0
		x"AB",x"F5",x"F4",x"7C",x"7A",x"3B",x"0D",x"8C", -- 0x00A8
		x"4B",x"55",x"BA",x"AA",x"5C",x"55",x"BB",x"AA", -- 0x00B0
		x"65",x"55",x"DA",x"AA",x"9D",x"54",x"34",x"AA", -- 0x00B8
		x"FD",x"7B",x"7E",x"27",x"C5",x"2B",x"0B",x"B5", -- 0x00C0
		x"FB",x"BD",x"7F",x"26",x"0F",x"1F",x"BF",x"EF", -- 0x00C8
		x"4B",x"51",x"B2",x"AB",x"7C",x"77",x"BB",x"AA", -- 0x00D0
		x"65",x"7D",x"DE",x"AA",x"99",x"94",x"D6",x"EA", -- 0x00D8
		x"ED",x"56",x"0D",x"0D",x"D7",x"AF",x"33",x"FF", -- 0x00E0
		x"4B",x"A6",x"F5",x"21",x"4B",x"0F",x"87",x"EF", -- 0x00E8
		x"CB",x"D7",x"BA",x"AA",x"DC",x"95",x"FB",x"EA", -- 0x00F0
		x"E5",x"F5",x"DA",x"AA",x"DD",x"F4",x"D4",x"EA", -- 0x00F8
		x"EC",x"44",x"11",x"51",x"F3",x"67",x"0B",x"3D", -- 0x0100
		x"5F",x"BD",x"7F",x"7F",x"5B",x"A3",x"E5",x"0C", -- 0x0108
		x"CB",x"D1",x"B2",x"AB",x"7C",x"F7",x"BB",x"AA", -- 0x0110
		x"65",x"7D",x"DE",x"AA",x"DB",x"56",x"B4",x"AA", -- 0x0118
		x"DF",x"AE",x"51",x"23",x"81",x"16",x"AF",x"F5", -- 0x0120
		x"E4",x"A2",x"50",x"B8",x"9C",x"9C",x"0C",x"6D", -- 0x0128
		x"CF",x"ED",x"5A",x"AA",x"FE",x"7D",x"7B",x"FA", -- 0x0130
		x"9D",x"CD",x"1E",x"1A",x"79",x"54",x"F4",x"EA", -- 0x0138
		x"FD",x"37",x"4B",x"37",x"41",x"03",x"0F",x"35", -- 0x0140
		x"EB",x"D5",x"97",x"CC",x"96",x"69",x"2B",x"D4", -- 0x0148
		x"CB",x"D5",x"96",x"AB",x"7C",x"77",x"BB",x"AA", -- 0x0150
		x"65",x"7D",x"DE",x"AA",x"99",x"74",x"14",x"AA", -- 0x0158
		x"FF",x"DD",x"DD",x"A9",x"90",x"EA",x"63",x"01", -- 0x0160
		x"88",x"F5",x"D3",x"C9",x"43",x"A0",x"98",x"FF", -- 0x0168
		x"CB",x"F1",x"FB",x"FF",x"FC",x"F8",x"C1",x"51", -- 0x0170
		x"4B",x"A3",x"8D",x"17",x"C7",x"0D",x"C1",x"F3", -- 0x0178
		x"55",x"AB",x"EA",x"D5",x"E5",x"EA",x"FA",x"FD", -- 0x0180
		x"FB",x"CD",x"14",x"7E",x"7E",x"9F",x"AF",x"4F", -- 0x0188
		x"4B",x"51",x"B2",x"AA",x"5C",x"55",x"BB",x"AA", -- 0x0190
		x"65",x"75",x"DA",x"AA",x"DB",x"F4",x"D4",x"EA", -- 0x0198
		x"EF",x"47",x"10",x"13",x"CB",x"7F",x"7E",x"B8", -- 0x01A0
		x"C3",x"0D",x"13",x"2C",x"D6",x"EB",x"25",x"D4", -- 0x01A8
		x"CF",x"0D",x"3A",x"EB",x"FC",x"F7",x"7B",x"EA", -- 0x01B0
		x"E5",x"7D",x"DE",x"AA",x"9D",x"56",x"54",x"AA", -- 0x01B8
		x"3F",x"DF",x"6C",x"F3",x"FA",x"AD",x"BB",x"D3", -- 0x01C0
		x"DF",x"E5",x"F1",x"4C",x"F2",x"EA",x"76",x"BC", -- 0x01C8
		x"F7",x"AB",x"DB",x"65",x"52",x"05",x"AE",x"DA", -- 0x01D0
		x"E3",x"47",x"06",x"0E",x"07",x"14",x"7C",x"EA", -- 0x01D8
		x"55",x"CB",x"3A",x"FF",x"BF",x"1F",x"5F",x"6E", -- 0x01E0
		x"AE",x"F8",x"6D",x"1E",x"4E",x"17",x"81",x"E3", -- 0x01E8
		x"4B",x"5D",x"BE",x"DF",x"7F",x"CF",x"8F",x"86", -- 0x01F0
		x"4B",x"55",x"E2",x"FB",x"67",x"19",x"14",x"FF", -- 0x01F8
		x"55",x"AB",x"AE",x"57",x"D6",x"EC",x"BD",x"31", -- 0x0200
		x"13",x"B9",x"5C",x"5E",x"68",x"96",x"AB",x"4F", -- 0x0208
		x"4B",x"5F",x"FF",x"FF",x"3F",x"DF",x"D7",x"CD", -- 0x0210
		x"AE",x"7D",x"B7",x"BF",x"9B",x"06",x"A9",x"CF", -- 0x0218
		x"55",x"AB",x"AA",x"55",x"D5",x"3A",x"52",x"D5", -- 0x0220
		x"2B",x"55",x"94",x"AD",x"B7",x"6D",x"2F",x"D7", -- 0x0228
		x"4B",x"51",x"B2",x"AA",x"5C",x"55",x"BB",x"AF", -- 0x0230
		x"6F",x"7E",x"FD",x"DA",x"8D",x"9F",x"09",x"1B", -- 0x0238
		x"57",x"AF",x"BF",x"59",x"F9",x"3D",x"5B",x"D0", -- 0x0240
		x"30",x"58",x"BF",x"BF",x"DF",x"77",x"30",x"F3", -- 0x0248
		x"C9",x"93",x"D5",x"E1",x"E2",x"63",x"5D",x"AB", -- 0x0250
		x"7F",x"37",x"37",x"9B",x"6A",x"B5",x"5F",x"27", -- 0x0258
		x"70",x"F2",x"E3",x"71",x"E7",x"CA",x"85",x"8C", -- 0x0260
		x"97",x"87",x"C9",x"C3",x"E7",x"62",x"31",x"F1", -- 0x0268
		x"5F",x"E7",x"AB",x"BF",x"DF",x"BD",x"17",x"6B", -- 0x0270
		x"FF",x"B7",x"37",x"9B",x"6A",x"75",x"DF",x"27", -- 0x0278
		x"60",x"B1",x"B1",x"58",x"E8",x"2C",x"54",x"D4", -- 0x0280
		x"2A",x"77",x"B5",x"EC",x"DA",x"7D",x"2D",x"C7", -- 0x0288
		x"DF",x"E7",x"6B",x"27",x"FF",x"7D",x"57",x"2B", -- 0x0290
		x"47",x"03",x"17",x"9B",x"8A",x"D5",x"DF",x"A7", -- 0x0298
		x"55",x"AB",x"BA",x"55",x"D5",x"2A",x"52",x"D5", -- 0x02A0
		x"2B",x"55",x"B6",x"ED",x"9A",x"69",x"25",x"D4", -- 0x02A8
		x"19",x"93",x"95",x"C1",x"42",x"63",x"B8",x"AE", -- 0x02B0
		x"67",x"55",x"DA",x"AA",x"DD",x"56",x"54",x"AA", -- 0x02B8
		x"FF",x"5E",x"17",x"96",x"C8",x"77",x"1F",x"06", -- 0x02C0
		x"CE",x"67",x"A3",x"F0",x"B0",x"6C",x"76",x"D5", -- 0x02C8
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"D7",x"EB", -- 0x02D0
		x"FF",x"77",x"77",x"DB",x"6A",x"55",x"5F",x"27", -- 0x02D8
		x"EE",x"47",x"17",x"11",x"DB",x"02",x"04",x"21", -- 0x02E0
		x"F0",x"D8",x"AF",x"C4",x"9A",x"69",x"25",x"D4", -- 0x02E8
		x"19",x"3E",x"2F",x"E5",x"43",x"E0",x"80",x"9C", -- 0x02F0
		x"2F",x"75",x"DA",x"AA",x"C9",x"26",x"54",x"AA", -- 0x02F8
		x"55",x"AB",x"AE",x"C7",x"F5",x"FA",x"B9",x"78", -- 0x0300
		x"9D",x"74",x"EF",x"36",x"70",x"29",x"BF",x"EF", -- 0x0308
		x"4B",x"55",x"B4",x"AB",x"F4",x"F3",x"FB",x"FF", -- 0x0310
		x"7C",x"F1",x"AE",x"CF",x"C7",x"69",x"34",x"FF", -- 0x0318
		x"55",x"AB",x"AA",x"55",x"D5",x"2B",x"57",x"DE", -- 0x0320
		x"F4",x"E6",x"6F",x"27",x"72",x"3B",x"9F",x"CF", -- 0x0328
		x"4B",x"51",x"B2",x"AA",x"54",x"FD",x"7F",x"7F", -- 0x0330
		x"FC",x"D9",x"E6",x"FB",x"A7",x"49",x"14",x"FF", -- 0x0338
		x"EE",x"47",x"15",x"56",x"E9",x"6C",x"05",x"03", -- 0x0340
		x"E1",x"D0",x"AF",x"AE",x"DA",x"6D",x"29",x"D4", -- 0x0348
		x"97",x"0B",x"1B",x"85",x"E2",x"D9",x"CF",x"C1", -- 0x0350
		x"C2",x"F1",x"D8",x"AC",x"9B",x"57",x"54",x"AA", -- 0x0358
		x"EF",x"52",x"19",x"03",x"85",x"C3",x"61",x"FE", -- 0x0360
		x"2F",x"55",x"97",x"AC",x"92",x"6D",x"29",x"D4", -- 0x0368
		x"E9",x"C6",x"EF",x"E3",x"45",x"E0",x"F0",x"AC", -- 0x0370
		x"67",x"7D",x"DE",x"AA",x"99",x"54",x"54",x"AA", -- 0x0378
		x"AE",x"6A",x"53",x"97",x"56",x"6E",x"A4",x"D4", -- 0x0380
		x"AE",x"AB",x"55",x"55",x"53",x"AB",x"AA",x"96", -- 0x0388
		x"1F",x"27",x"2B",x"1F",x"17",x"2D",x"17",x"6B", -- 0x0390
		x"3B",x"17",x"35",x"1B",x"6A",x"35",x"1F",x"27", -- 0x0398
		x"AF",x"5F",x"5F",x"BF",x"27",x"D3",x"8B",x"90", -- 0x03A0
		x"80",x"C0",x"42",x"40",x"62",x"97",x"BC",x"2B", -- 0x03A8
		x"94",x"E6",x"E9",x"FC",x"FF",x"FE",x"FE",x"FF", -- 0x03B0
		x"3E",x"0E",x"4D",x"35",x"52",x"C9",x"A7",x"55", -- 0x03B8
		x"AA",x"D4",x"D1",x"E2",x"07",x"DB",x"8B",x"31", -- 0x03C0
		x"91",x"88",x"08",x"45",x"63",x"88",x"D4",x"2B", -- 0x03C8
		x"B4",x"4A",x"55",x"35",x"89",x"CA",x"E0",x"E1", -- 0x03D0
		x"72",x"F2",x"E5",x"C5",x"02",x"29",x"AB",x"55", -- 0x03D8
		x"4C",x"16",x"23",x"AF",x"59",x"5A",x"10",x"90", -- 0x03E0
		x"68",x"29",x"D4",x"57",x"2C",x"AA",x"44",x"36", -- 0x03E8
		x"0A",x"D4",x"E3",x"F8",x"FA",x"FB",x"BD",x"7C", -- 0x03F0
		x"5E",x"3C",x"19",x"3A",x"D2",x"15",x"C8",x"26", -- 0x03F8
		x"07",x"01",x"03",x"01",x"01",x"00",x"00",x"00", -- 0x0400
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0408
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"5F",x"2F", -- 0x0410
		x"1F",x"05",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x0418
		x"FF",x"7F",x"1F",x"1F",x"07",x"03",x"07",x"03", -- 0x0420
		x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0428
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0430
		x"FF",x"FF",x"FD",x"5C",x"30",x"00",x"00",x"00", -- 0x0438
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"BF", -- 0x0440
		x"2F",x"1F",x"07",x"03",x"00",x"00",x"00",x"00", -- 0x0448
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0450
		x"FF",x"FF",x"FB",x"6C",x"A0",x"80",x"00",x"00", -- 0x0458
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0460
		x"FF",x"FF",x"BF",x"1F",x"25",x"00",x"00",x"00", -- 0x0468
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0470
		x"FF",x"FE",x"FF",x"B4",x"F0",x"80",x"00",x"00", -- 0x0478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0480
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"3F",x"00", -- 0x0488
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0490
		x"FF",x"FE",x"FB",x"F4",x"F0",x"C0",x"40",x"00", -- 0x0498
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"80", -- 0x04A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04B0
		x"FF",x"FF",x"FA",x"FC",x"F0",x"C0",x"00",x"00", -- 0x04B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FD", -- 0x04C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04D0
		x"FF",x"FF",x"FD",x"EC",x"E0",x"80",x"00",x"00", -- 0x04D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04F0
		x"FF",x"FF",x"FA",x"FC",x"F0",x"D0",x"E0",x"E0", -- 0x04F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"DF", -- 0x0500
		x"3F",x"0B",x"06",x"00",x"00",x"00",x"00",x"00", -- 0x0508
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FB", -- 0x0510
		x"DC",x"70",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x0518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0520
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"1F",x"00", -- 0x0528
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FD", -- 0x0530
		x"F4",x"F8",x"F0",x"D0",x"C0",x"80",x"40",x"00", -- 0x0538
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0540
		x"FF",x"FF",x"FE",x"FA",x"F4",x"E0",x"C0",x"80", -- 0x0548
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF", -- 0x0550
		x"EC",x"E0",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x0558
		x"FF",x"7F",x"3F",x"0B",x"07",x"01",x"01",x"00", -- 0x0560
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0568
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x0570
		x"FF",x"7F",x"7F",x"3F",x"3F",x"16",x"0C",x"00", -- 0x0578
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0580
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"17",x"00", -- 0x0588
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0590
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"F8",x"00", -- 0x0598
		x"00",x"00",x"01",x"00",x"01",x"03",x"02",x"01", -- 0x05A0
		x"03",x"03",x"02",x"00",x"01",x"01",x"00",x"00", -- 0x05A8
		x"7F",x"3F",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05B0
		x"7F",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"FF", -- 0x05B8
		x"07",x"03",x"0F",x"0B",x"0F",x"1F",x"0F",x"1F", -- 0x05C0
		x"17",x"0F",x"1F",x"07",x"0F",x"0B",x"07",x"07", -- 0x05C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05D8
		x"3F",x"3F",x"7F",x"5F",x"7F",x"7F",x"7F",x"7F", -- 0x05E0
		x"7F",x"7F",x"7F",x"7F",x"3F",x"7F",x"1F",x"3F", -- 0x05E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F8
		x"00",x"00",x"01",x"01",x"00",x"01",x"00",x"00", -- 0x0600
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0608
		x"7F",x"DF",x"FF",x"7F",x"FF",x"FF",x"FF",x"BF", -- 0x0610
		x"7F",x"5F",x"4F",x"1F",x"07",x"07",x"07",x"01", -- 0x0618
		x"05",x"07",x"0F",x"07",x"3F",x"17",x"0F",x"1F", -- 0x0620
		x"05",x"02",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x0628
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0630
		x"FF",x"FF",x"FF",x"3F",x"0F",x"07",x"07",x"01", -- 0x0638
		x"3F",x"3F",x"3F",x"3F",x"3F",x"1F",x"1F",x"1F", -- 0x0640
		x"07",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0650
		x"FF",x"FF",x"7F",x"1F",x"0F",x"07",x"07",x"01", -- 0x0658
		x"FF",x"7F",x"3F",x"3F",x"3F",x"1F",x"0F",x"1F", -- 0x0660
		x"17",x"0F",x"0F",x"05",x"03",x"00",x"00",x"00", -- 0x0668
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"47",x"01", -- 0x0678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0680
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FD", -- 0x0688
		x"FF",x"FE",x"FC",x"FC",x"FC",x"F8",x"F8",x"FC", -- 0x0690
		x"F8",x"F0",x"F0",x"E0",x"C0",x"80",x"00",x"00", -- 0x0698
		x"3F",x"5F",x"3F",x"7F",x"7F",x"3F",x"1F",x"1F", -- 0x06A0
		x"07",x"05",x"03",x"01",x"01",x"00",x"01",x"00", -- 0x06A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06B0
		x"FF",x"FF",x"FF",x"7F",x"FF",x"7F",x"BF",x"FF", -- 0x06B8
		x"05",x"07",x"0B",x"0F",x"37",x"17",x"0F",x"0F", -- 0x06C0
		x"0B",x"07",x"02",x"00",x"01",x"00",x"01",x"00", -- 0x06C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06D0
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"BF",x"FF", -- 0x06D8
		x"07",x"03",x"0F",x"07",x"0F",x"1F",x"0F",x"3F", -- 0x06E0
		x"5F",x"7F",x"7F",x"7F",x"3F",x"7F",x"3F",x"3F", -- 0x06E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0700
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0708
		x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"FC", -- 0x0710
		x"FC",x"F8",x"F8",x"F8",x"E0",x"F0",x"A0",x"E0", -- 0x0718
		x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"1C", -- 0x0720
		x"0C",x"2E",x"0A",x"34",x"11",x"07",x"3A",x"0E", -- 0x0728
		x"BF",x"3F",x"5F",x"3F",x"2F",x"19",x"07",x"66", -- 0x0730
		x"37",x"7B",x"F9",x"5B",x"62",x"BD",x"4B",x"A7", -- 0x0738
		x"2B",x"67",x"15",x"2A",x"26",x"09",x"1C",x"08", -- 0x0740
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0748
		x"F7",x"AB",x"7B",x"B7",x"52",x"05",x"2F",x"1E", -- 0x0750
		x"0B",x"17",x"03",x"00",x"21",x"1B",x"3F",x"FF", -- 0x0758
		x"2E",x"DF",x"56",x"0A",x"D0",x"60",x"60",x"20", -- 0x0760
		x"D0",x"38",x"18",x"00",x"08",x"94",x"FC",x"FD", -- 0x0768
		x"B8",x"2E",x"12",x"00",x"00",x"00",x"00",x"00", -- 0x0770
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
		x"55",x"AB",x"AE",x"57",x"D5",x"2B",x"53",x"D5", -- 0x0780
		x"2B",x"55",x"B7",x"AC",x"D2",x"6D",x"25",x"D4", -- 0x0788
		x"4B",x"55",x"B6",x"AB",x"7C",x"77",x"BB",x"AA", -- 0x0790
		x"65",x"7D",x"DE",x"AA",x"DB",x"56",x"55",x"AA", -- 0x0798
		x"55",x"AB",x"AA",x"55",x"D5",x"2A",x"52",x"D5", -- 0x07A0
		x"2B",x"55",x"D6",x"AD",x"92",x"65",x"29",x"D6", -- 0x07A8
		x"4B",x"55",x"B6",x"AA",x"5C",x"55",x"BB",x"AA", -- 0x07B0
		x"65",x"75",x"DA",x"AA",x"9B",x"56",x"34",x"AA", -- 0x07B8
		x"B3",x"D5",x"E6",x"4A",x"AD",x"B6",x"D8",x"65", -- 0x07C0
		x"95",x"EA",x"6D",x"96",x"D9",x"66",x"9B",x"CD", -- 0x07C8
		x"B5",x"5B",x"64",x"B7",x"45",x"9A",x"EC",x"6B", -- 0x07D0
		x"96",x"A9",x"2E",x"D5",x"29",x"EA",x"17",x"D9", -- 0x07D8
		x"55",x"AA",x"19",x"B5",x"52",x"49",x"A7",x"9A", -- 0x07E0
		x"6A",x"95",x"D2",x"69",x"A6",x"99",x"6C",x"B6", -- 0x07E8
		x"5A",x"A5",x"9B",x"48",x"BA",x"65",x"13",x"96", -- 0x07F0
		x"69",x"56",x"D1",x"2A",x"D6",x"15",x"E9",x"A6", -- 0x07F8
		x"00",x"EF",x"DF",x"A6",x"60",x"00",x"00",x"7F", -- 0x0800
		x"7F",x"7F",x"7F",x"03",x"03",x"03",x"03",x"03", -- 0x0808
		x"00",x"FE",x"FE",x"56",x"2E",x"0E",x"16",x"8E", -- 0x0810
		x"8E",x"8E",x"8E",x"86",x"B6",x"8E",x"8E",x"8E", -- 0x0818
		x"03",x"03",x"03",x"03",x"03",x"00",x"00",x"00", -- 0x0820
		x"00",x"00",x"01",x"26",x"8B",x"C7",x"FF",x"FF", -- 0x0828
		x"9E",x"86",x"8C",x"BA",x"BE",x"2E",x"1A",x"3E", -- 0x0830
		x"1E",x"9E",x"5E",x"BE",x"FE",x"2E",x"1E",x"9E", -- 0x0838
		x"FF",x"8B",x"C1",x"F3",x"FF",x"3E",x"0F",x"03", -- 0x0840
		x"E7",x"BF",x"2F",x"9F",x"8F",x"C3",x"E7",x"E3", -- 0x0848
		x"0E",x"BE",x"B6",x"BE",x"6E",x"1E",x"7E",x"F6", -- 0x0850
		x"DE",x"9E",x"AE",x"0E",x"1E",x"16",x"AE",x"BE", -- 0x0858
		x"EF",x"77",x"67",x"C2",x"E0",x"F2",x"B7",x"9F", -- 0x0860
		x"F9",x"F3",x"39",x"18",x"08",x"4E",x"00",x"00", -- 0x0868
		x"16",x"8E",x"9E",x"7E",x"7E",x"FE",x"BE",x"2E", -- 0x0870
		x"9E",x"9E",x"2E",x"7E",x"3E",x"3E",x"00",x"00", -- 0x0878
		x"00",x"1E",x"F7",x"B4",x"38",x"56",x"EF",x"F6", -- 0x0880
		x"EE",x"A7",x"03",x"82",x"E1",x"E5",x"C6",x"86", -- 0x0888
		x"00",x"68",x"28",x"3C",x"5C",x"3E",x"D4",x"EA", -- 0x0890
		x"FE",x"76",x"76",x"FA",x"68",x"D8",x"EC",x"F8", -- 0x0898
		x"DF",x"8D",x"C5",x"C4",x"E0",x"E2",x"C7",x"EF", -- 0x08A0
		x"EF",x"C7",x"87",x"01",x"43",x"70",x"79",x"BF", -- 0x08A8
		x"EC",x"7C",x"3E",x"2E",x"10",x"04",x"0C",x"FA", -- 0x08B0
		x"FC",x"7E",x"3C",x"DC",x"56",x"E6",x"E4",x"F0", -- 0x08B8
		x"DF",x"3E",x"37",x"04",x"80",x"CE",x"FF",x"76", -- 0x08C0
		x"6E",x"27",x"43",x"02",x"41",x"E5",x"F6",x"CE", -- 0x08C8
		x"5C",x"64",x"06",x"1C",x"58",x"3E",x"DC",x"EE", -- 0x08D0
		x"FE",x"76",x"60",x"D4",x"6C",x"DE",x"DE",x"E6", -- 0x08D8
		x"9F",x"85",x"C1",x"CC",x"70",x"22",x"77",x"3F", -- 0x08E0
		x"0E",x"07",x"87",x"E0",x"F3",x"24",x"00",x"00", -- 0x08E8
		x"EE",x"5E",x"1C",x"2A",x"04",x"8C",x"FE",x"FE", -- 0x08F0
		x"FC",x"DE",x"3E",x"12",x"0C",x"88",x"00",x"00", -- 0x08F8
		x"00",x"3F",x"27",x"0F",x"07",x"2A",x"0C",x"28", -- 0x0900
		x"3C",x"0C",x"1E",x"0E",x"1E",x"04",x"3C",x"00", -- 0x0908
		x"00",x"FF",x"FF",x"57",x"04",x"80",x"00",x"7C", -- 0x0910
		x"7C",x"7C",x"7C",x"00",x"00",x"00",x"00",x"00", -- 0x0918
		x"1E",x"0F",x"32",x"3A",x"0C",x"3E",x"1D",x"1E", -- 0x0920
		x"3E",x"0B",x"07",x"3E",x"0F",x"07",x"2F",x"0B", -- 0x0928
		x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00", -- 0x0930
		x"00",x"04",x"4C",x"A6",x"16",x"82",x"C5",x"E7", -- 0x0938
		x"07",x"21",x"33",x"3E",x"3E",x"1C",x"0C",x"1E", -- 0x0940
		x"0E",x"1C",x"0B",x"0F",x"07",x"0B",x"02",x"01", -- 0x0948
		x"EB",x"E7",x"F0",x"7A",x"DF",x"7F",x"2B",x"31", -- 0x0950
		x"7F",x"6F",x"FF",x"97",x"8F",x"C3",x"E3",x"F3", -- 0x0958
		x"37",x"25",x"32",x"15",x"0B",x"09",x"05",x"04", -- 0x0960
		x"22",x"31",x"3A",x"21",x"20",x"31",x"00",x"00", -- 0x0968
		x"FC",x"BD",x"1E",x"77",x"EF",x"A2",x"71",x"99", -- 0x0970
		x"0F",x"85",x"9B",x"02",x"80",x"C1",x"00",x"00", -- 0x0978
		x"00",x"03",x"17",x"24",x"20",x"16",x"3F",x"16", -- 0x0980
		x"0E",x"0F",x"07",x"02",x"00",x"1A",x"1E",x"2F", -- 0x0988
		x"00",x"F7",x"EB",x"DF",x"4F",x"05",x"C5",x"EB", -- 0x0990
		x"FF",x"77",x"75",x"F0",x"D9",x"4F",x"4F",x"FF", -- 0x0998
		x"17",x"2F",x"0B",x"07",x"03",x"01",x"03",x"3B", -- 0x09A0
		x"11",x"12",x"37",x"03",x"27",x"1F",x"07",x"2F", -- 0x09A8
		x"EF",x"FF",x"FF",x"F7",x"BF",x"FD",x"FF",x"FF", -- 0x09B0
		x"FF",x"7F",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE", -- 0x09B8
		x"07",x"03",x"03",x"37",x"1F",x"1B",x"27",x"27", -- 0x09C0
		x"07",x"03",x"03",x"2F",x"13",x"11",x"37",x"07", -- 0x09C8
		x"F4",x"FC",x"FC",x"FE",x"DF",x"EF",x"FE",x"FC", -- 0x09D0
		x"FC",x"FC",x"FE",x"DE",x"FF",x"FF",x"FF",x"FF", -- 0x09D8
		x"07",x"13",x"3F",x"25",x"03",x"01",x"3B",x"1F", -- 0x09E0
		x"1F",x"1F",x"3F",x"3F",x"17",x"0C",x"00",x"00", -- 0x09E8
		x"FD",x"FB",x"FF",x"FF",x"FF",x"BE",x"FE",x"F6", -- 0x09F0
		x"EF",x"C5",x"C1",x"F7",x"BD",x"51",x"00",x"00", -- 0x09F8
		x"FF",x"FF",x"E0",x"C0",x"C0",x"C0",x"F1",x"E1", -- 0x0A00
		x"C1",x"C1",x"C3",x"C7",x"E3",x"C3",x"C3",x"C3", -- 0x0A08
		x"FF",x"FF",x"7F",x"7E",x"7C",x"F8",x"F0",x"F0", -- 0x0A10
		x"E0",x"E0",x"C0",x"C0",x"81",x"81",x"83",x"83", -- 0x0A18
		x"C7",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC", -- 0x0A20
		x"FC",x"FC",x"FC",x"F8",x"F8",x"FF",x"FF",x"F8", -- 0x0A28
		x"07",x"07",x"0F",x"08",x"00",x"00",x"00",x"10", -- 0x0A30
		x"11",x"13",x"03",x"03",x"07",x"FF",x"FF",x"3F", -- 0x0A38
		x"F0",x"F0",x"F0",x"F0",x"F0",x"E0",x"E0",x"E0", -- 0x0A40
		x"E0",x"C0",x"C0",x"C1",x"C1",x"81",x"83",x"83", -- 0x0A48
		x"31",x"61",x"61",x"61",x"63",x"71",x"E1",x"E1", -- 0x0A50
		x"E1",x"E1",x"E1",x"E1",x"E1",x"E1",x"E3",x"E3", -- 0x0A58
		x"03",x"07",x"07",x"07",x"0F",x"1F",x"3C",x"38", -- 0x0A60
		x"78",x"60",x"C0",x"C0",x"C0",x"C0",x"FF",x"FF", -- 0x0A68
		x"C3",x"C7",x"FF",x"FF",x"E1",x"C1",x"01",x"01", -- 0x0A70
		x"01",x"01",x"81",x"01",x"03",x"07",x"FF",x"FF", -- 0x0A78
		x"FF",x"FF",x"DF",x"DF",x"C3",x"FF",x"FF",x"EF", -- 0x0A80
		x"CF",x"CF",x"C0",x"C1",x"FD",x"DD",x"DD",x"C4", -- 0x0A88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"DF",x"DF", -- 0x0A90
		x"DF",x"C3",x"FF",x"EF",x"EF",x"EF",x"E3",x"7F", -- 0x0A98
		x"E1",x"C0",x"C2",x"FE",x"EE",x"CF",x"CE",x"C2", -- 0x0AA0
		x"C6",x"FF",x"FF",x"FF",x"EF",x"CE",x"CE",x"C3", -- 0x0AA8
		x"FF",x"F7",x"F7",x"F7",x"13",x"E1",x"C1",x"C1", -- 0x0AB0
		x"43",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"CF", -- 0x0AB8
		x"C7",x"FF",x"DD",x"DD",x"DD",x"DC",x"C7",x"FE", -- 0x0AC0
		x"FE",x"FF",x"FF",x"FF",x"DF",x"DE",x"DE",x"DE", -- 0x0AC8
		x"C3",x"F7",x"FF",x"FF",x"F7",x"17",x"F7",x"F7", -- 0x0AD0
		x"37",x"F3",x"FF",x"DF",x"1F",x"1F",x"1F",x"1F", -- 0x0AD8
		x"DE",x"C2",x"FF",x"FF",x"EF",x"CF",x"CF",x"CF", -- 0x0AE0
		x"C0",x"C1",x"FF",x"F7",x"F7",x"F0",x"FF",x"FF", -- 0x0AE8
		x"03",x"7F",x"BF",x"BF",x"87",x"E1",x"C1",x"C3", -- 0x0AF0
		x"FF",x"DF",x"DF",x"DF",x"DF",x"C3",x"FF",x"FF", -- 0x0AF8
		x"FF",x"F8",x"B0",x"B1",x"B8",x"B0",x"B0",x"91", -- 0x0B00
		x"FF",x"FF",x"FF",x"FF",x"DE",x"DC",x"DC",x"DC", -- 0x0B08
		x"FF",x"FF",x"BF",x"3F",x"3F",x"3F",x"03",x"07", -- 0x0B10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B18
		x"C4",x"FE",x"EF",x"CE",x"CE",x"CE",x"C2",x"C6", -- 0x0B20
		x"FF",x"EF",x"CF",x"CF",x"CF",x"C1",x"C3",x"FF", -- 0x0B28
		x"03",x"1F",x"1F",x"1F",x"03",x"21",x"01",x"43", -- 0x0B30
		x"FF",x"BF",x"3F",x"3F",x"3F",x"03",x"07",x"FF", -- 0x0B38
		x"EF",x"CF",x"CC",x"CD",x"CE",x"CC",x"CC",x"CC", -- 0x0B40
		x"C7",x"CF",x"FF",x"FF",x"FF",x"EF",x"CF",x"C1", -- 0x0B48
		x"BF",x"BF",x"3F",x"3F",x"3F",x"3F",x"03",x"07", -- 0x0B50
		x"FF",x"FF",x"FF",x"8F",x"0F",x"0F",x"0F",x"2F", -- 0x0B58
		x"C3",x"FF",x"DF",x"DF",x"DF",x"C1",x"FF",x"EF", -- 0x0B60
		x"CF",x"CF",x"CF",x"CF",x"C0",x"C1",x"FF",x"FF", -- 0x0B68
		x"E3",x"71",x"61",x"61",x"63",x"3F",x"DF",x"9F", -- 0x0B70
		x"9F",x"9F",x"9F",x"9F",x"83",x"87",x"FF",x"FF", -- 0x0B78
		x"FF",x"FF",x"E1",x"C1",x"C0",x"C0",x"C1",x"C1", -- 0x0B80
		x"C3",x"E0",x"C0",x"C0",x"C0",x"C1",x"FF",x"FF", -- 0x0B88
		x"FF",x"DF",x"FF",x"7F",x"3F",x"1F",x"97",x"87", -- 0x0B90
		x"DF",x"9F",x"8F",x"E7",x"BF",x"0F",x"27",x"FF", -- 0x0B98
		x"FF",x"FC",x"D8",x"D8",x"D8",x"D8",x"D8",x"C0", -- 0x0BA0
		x"FF",x"DF",x"DE",x"DE",x"C3",x"FE",x"DE",x"DE", -- 0x0BA8
		x"FF",x"FF",x"BF",x"3F",x"3F",x"3F",x"3F",x"03", -- 0x0BB0
		x"07",x"3F",x"1F",x"5F",x"DF",x"DF",x"DF",x"DF", -- 0x0BB8
		x"DE",x"C6",x"FF",x"EF",x"CF",x"CF",x"CF",x"C1", -- 0x0BC0
		x"C3",x"FF",x"FF",x"FF",x"EF",x"CE",x"CE",x"C2", -- 0x0BC8
		x"C3",x"79",x"F1",x"71",x"71",x"71",x"73",x"1F", -- 0x0BD0
		x"FF",x"FF",x"FF",x"EF",x"EF",x"EF",x"E3",x"FF", -- 0x0BD8
		x"C6",x"E0",x"C1",x"C1",x"C0",x"C2",x"FF",x"EF", -- 0x0BE0
		x"CF",x"CF",x"CF",x"CF",x"C0",x"C1",x"FF",x"FF", -- 0x0BE8
		x"FF",x"2F",x"EF",x"0F",x"0F",x"23",x"FF",x"FF", -- 0x0BF0
		x"DF",x"9F",x"9F",x"9F",x"83",x"87",x"FF",x"FF", -- 0x0BF8
		x"FF",x"FF",x"FB",x"FB",x"FB",x"F8",x"FF",x"DE", -- 0x0C00
		x"DE",x"DE",x"DF",x"C2",x"FE",x"BE",x"83",x"FF", -- 0x0C08
		x"FF",x"FF",x"EF",x"CF",x"CF",x"43",x"07",x"3F", -- 0x0C10
		x"1F",x"5F",x"03",x"3F",x"1F",x"43",x"FF",x"7F", -- 0x0C18
		x"DB",x"C9",x"FF",x"FF",x"FF",x"BB",x"B3",x"B3", -- 0x0C20
		x"93",x"F3",x"B0",x"B1",x"BF",x"9F",x"FF",x"FF", -- 0x0C28
		x"7F",x"7F",x"07",x"FF",x"FF",x"BF",x"BF",x"BF", -- 0x0C30
		x"87",x"87",x"E7",x"67",x"63",x"67",x"3F",x"FF", -- 0x0C38
		x"FF",x"FF",x"FD",x"FD",x"FC",x"07",x"E1",x"C0", -- 0x0C40
		x"C0",x"C0",x"C3",x"7F",x"FF",x"FF",x"FF",x"EF", -- 0x0C48
		x"FF",x"FF",x"F9",x"F1",x"11",x"FB",x"7F",x"7F", -- 0x0C50
		x"0F",x"1F",x"FF",x"FF",x"F3",x"63",x"63",x"67", -- 0x0C58
		x"EF",x"EF",x"E1",x"FE",x"1C",x"C4",x"FF",x"7B", -- 0x0C60
		x"73",x"33",x"F3",x"F3",x"F0",x"30",x"FF",x"FF", -- 0x0C68
		x"3F",x"DF",x"DF",x"1F",x"1F",x"43",x"FF",x"F7", -- 0x0C70
		x"F3",x"F1",x"E1",x"E1",x"61",x"E3",x"FF",x"FF", -- 0x0C78
		x"FF",x"F7",x"FD",x"FF",x"FF",x"FF",x"3F",x"76", -- 0x0C80
		x"FE",x"FF",x"7D",x"6D",x"7D",x"FC",x"FF",x"FF", -- 0x0C88
		x"FF",x"F9",x"71",x"71",x"71",x"03",x"11",x"01", -- 0x0C90
		x"23",x"FF",x"BF",x"BF",x"BF",x"83",x"FF",x"FF", -- 0x0C98
		x"FF",x"F8",x"F0",x"F1",x"FF",x"17",x"E7",x"E7", -- 0x0CA0
		x"E7",x"E0",x"E1",x"F8",x"30",x"70",x"FF",x"FF", -- 0x0CA8
		x"FF",x"FF",x"BF",x"BF",x"BF",x"83",x"FF",x"DF", -- 0x0CB0
		x"DF",x"DF",x"DF",x"47",x"7F",x"FF",x"FF",x"FF", -- 0x0CB8
		x"FF",x"FF",x"31",x"21",x"21",x"21",x"23",x"3F", -- 0x0CC0
		x"3E",x"9F",x"1F",x"33",x"17",x"03",x"84",x"F0", -- 0x0CC8
		x"FF",x"FF",x"FF",x"DF",x"3F",x"2F",x"27",x"1F", -- 0x0CD0
		x"4F",x"1F",x"8B",x"C3",x"C7",x"7F",x"7F",x"FF", -- 0x0CD8
		x"FF",x"FF",x"EF",x"EF",x"EF",x"E0",x"FF",x"2E", -- 0x0CE0
		x"EE",x"EF",x"E2",x"FE",x"DE",x"42",x"FF",x"FF", -- 0x0CE8
		x"FF",x"FF",x"BF",x"BF",x"BF",x"83",x"F1",x"E1", -- 0x0CF0
		x"23",x"3F",x"1F",x"1F",x"1F",x"43",x"FF",x"FF", -- 0x0CF8
		x"FF",x"FF",x"EF",x"CF",x"CF",x"CF",x"C0",x"C0", -- 0x0D00
		x"FF",x"FF",x"FF",x"DF",x"DE",x"DE",x"DE",x"C2", -- 0x0D08
		x"FF",x"FF",x"EF",x"CF",x"FF",x"FF",x"00",x"01", -- 0x0D10
		x"FF",x"FF",x"FF",x"07",x"07",x"07",x"07",x"17", -- 0x0D18
		x"FF",x"DD",x"DD",x"DD",x"DC",x"C7",x"FE",x"DC", -- 0x0D20
		x"DC",x"C4",x"FC",x"DC",x"DC",x"C4",x"FF",x"FF", -- 0x0D28
		x"F1",x"FF",x"FF",x"EF",x"2F",x"EF",x"EF",x"EF", -- 0x0D30
		x"E1",x"FF",x"EF",x"E1",x"3F",x"6F",x"E3",x"FF", -- 0x0D38
		x"FF",x"FF",x"DF",x"DF",x"DF",x"C1",x"FF",x"DF", -- 0x0D40
		x"DE",x"DE",x"C3",x"E0",x"C0",x"C0",x"C0",x"C3", -- 0x0D48
		x"FF",x"FF",x"BF",x"3E",x"3E",x"06",x"0F",x"0F", -- 0x0D50
		x"07",x"17",x"F7",x"F0",x"FF",x"FF",x"1F",x"FF", -- 0x0D58
		x"FF",x"FF",x"FD",x"F9",x"F9",x"F8",x"D8",x"DE", -- 0x0D60
		x"DC",x"DC",x"DF",x"DE",x"DE",x"C2",x"FE",x"FF", -- 0x0D68
		x"FF",x"FB",x"FB",x"FB",x"F8",x"1C",x"38",x"18", -- 0x0D70
		x"18",x"39",x"0F",x"0B",x"0B",x"08",x"1F",x"FF", -- 0x0D78
		x"FF",x"FF",x"EF",x"EF",x"EF",x"E0",x"FC",x"D8", -- 0x0D80
		x"D8",x"D8",x"D8",x"DE",x"DC",x"C4",x"FF",x"FF", -- 0x0D88
		x"FF",x"EF",x"FF",x"F7",x"E7",x"E7",x"60",x"60", -- 0x0D90
		x"7F",x"7F",x"F8",x"70",x"70",x"F0",x"FF",x"FF", -- 0x0D98
		x"FF",x"E3",x"C3",x"C5",x"FD",x"DD",x"DD",x"DD", -- 0x0DA0
		x"C4",x"F1",x"E0",x"E2",x"FE",x"DE",x"C3",x"FF", -- 0x0DA8
		x"FF",x"FF",x"FE",x"F6",x"F6",x"F6",x"F3",x"FF", -- 0x0DB0
		x"3B",x"F3",x"F3",x"F3",x"F0",x"30",x"FF",x"FF", -- 0x0DB8
		x"FF",x"E0",x"C0",x"C1",x"FF",x"DF",x"C7",x"E5", -- 0x0DC0
		x"C1",x"C1",x"C9",x"F9",x"D8",x"C8",x"FF",x"FF", -- 0x0DC8
		x"FF",x"FF",x"7F",x"7E",x"7E",x"06",x"FE",x"FE", -- 0x0DD0
		x"FE",x"DF",x"DF",x"DF",x"43",x"FF",x"FF",x"FF", -- 0x0DD8
		x"FF",x"FF",x"DF",x"DC",x"D8",x"D8",x"C8",x"E0", -- 0x0DE0
		x"C0",x"CF",x"F7",x"E7",x"E0",x"E0",x"FF",x"FF", -- 0x0DE8
		x"FF",x"F3",x"E3",x"61",x"65",x"7D",x"7D",x"7C", -- 0x0DF0
		x"FF",x"FE",x"FE",x"FE",x"1E",x"3E",x"FF",x"FF", -- 0x0DF8
		x"FF",x"FF",x"FD",x"D9",x"D8",x"D8",x"DF",x"CB", -- 0x0E00
		x"F9",x"FF",x"F3",x"E1",x"E1",x"E1",x"E4",x"FF", -- 0x0E08
		x"FF",x"F9",x"F1",x"F1",x"11",x"33",x"FF",x"7F", -- 0x0E10
		x"07",x"FF",x"FF",x"FF",x"F7",x"F7",x"17",x"F7", -- 0x0E18
		x"FE",x"FE",x"FE",x"9F",x"9B",x"8F",x"87",x"CF", -- 0x0E20
		x"C2",x"F0",x"F9",x"F9",x"F8",x"F8",x"FE",x"FF", -- 0x0E28
		x"03",x"09",x"11",x"F1",x"F1",x"F3",x"FF",x"FF", -- 0x0E30
		x"FF",x"FF",x"FF",x"7F",x"AF",x"4F",x"2F",x"FF", -- 0x0E38
		x"FF",x"FF",x"FF",x"BF",x"3F",x"3F",x"3F",x"06", -- 0x0E40
		x"0E",x"FE",x"FE",x"FF",x"5F",x"1F",x"1F",x"9F", -- 0x0E48
		x"FF",x"FF",x"7F",x"7F",x"7F",x"07",x"3F",x"1F", -- 0x0E50
		x"1F",x"1F",x"5F",x"C3",x"FF",x"FF",x"FF",x"7F", -- 0x0E58
		x"1F",x"07",x"0F",x"FE",x"EE",x"EE",x"EF",x"E6", -- 0x0E60
		x"3E",x"FE",x"7E",x"7E",x"7E",x"07",x"FF",x"FF", -- 0x0E68
		x"7F",x"07",x"3F",x"1F",x"1F",x"5F",x"C3",x"FF", -- 0x0E70
		x"DF",x"DF",x"DF",x"DF",x"5F",x"C7",x"FF",x"FF", -- 0x0E78
		x"FF",x"FF",x"DD",x"D9",x"D9",x"D9",x"C9",x"F8", -- 0x0E80
		x"FF",x"EF",x"CF",x"CF",x"CF",x"C1",x"C3",x"E2", -- 0x0E88
		x"FF",x"FF",x"FF",x"87",x"87",x"E7",x"E7",x"E3", -- 0x0E90
		x"E7",x"FF",x"BF",x"BF",x"87",x"FF",x"FF",x"EF", -- 0x0E98
		x"C0",x"C0",x"C0",x"C4",x"FC",x"FC",x"DC",x"DF", -- 0x0EA0
		x"DF",x"DF",x"DF",x"DF",x"C0",x"FF",x"FF",x"FF", -- 0x0EA8
		x"EF",x"EF",x"E3",x"F3",x"E3",x"23",x"67",x"FF", -- 0x0EB0
		x"FF",x"DF",x"DF",x"DF",x"43",x"FF",x"FF",x"FF", -- 0x0EB8
		x"FF",x"FF",x"DF",x"DF",x"C0",x"FE",x"DE",x"DC", -- 0x0EC0
		x"DC",x"C4",x"FF",x"F7",x"F7",x"F7",x"F0",x"FF", -- 0x0EC8
		x"FF",x"FF",x"7F",x"7F",x"07",x"07",x"07",x"07", -- 0x0ED0
		x"03",x"1F",x"DF",x"DF",x"9F",x"9F",x"07",x"8F", -- 0x0ED8
		x"FF",x"FD",x"B9",x"B9",x"B9",x"B9",x"B8",x"98", -- 0x0EE0
		x"FF",x"DE",x"C2",x"E0",x"C0",x"C2",x"FF",x"FF", -- 0x0EE8
		x"FF",x"F9",x"F1",x"F1",x"F1",x"F1",x"13",x"3F", -- 0x0EF0
		x"FF",x"DF",x"DF",x"DF",x"DF",x"43",x"FF",x"FF", -- 0x0EF8
		x"FF",x"FF",x"DE",x"C2",x"FE",x"DF",x"DF",x"DF", -- 0x0F00
		x"DF",x"C3",x"FF",x"FF",x"FF",x"F0",x"E0",x"E0", -- 0x0F08
		x"FF",x"1F",x"0F",x"0F",x"21",x"FF",x"BF",x"3F", -- 0x0F10
		x"01",x"03",x"FF",x"FF",x"FF",x"5F",x"5F",x"47", -- 0x0F18
		x"E0",x"FF",x"FF",x"EE",x"CE",x"CE",x"CF",x"CE", -- 0x0F20
		x"CE",x"CF",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF", -- 0x0F28
		x"F7",x"B7",x"F7",x"F7",x"F1",x"18",x"00",x"00", -- 0x0F30
		x"10",x"F0",x"F1",x"FF",x"17",x"31",x"FF",x"FF", -- 0x0F38
		x"FF",x"FB",x"EF",x"E7",x"9F",x"8B",x"87",x"C1", -- 0x0F40
		x"F3",x"FF",x"FF",x"E1",x"C1",x"C0",x"C0",x"C2", -- 0x0F48
		x"FF",x"F0",x"E0",x"E0",x"E0",x"E1",x"E3",x"C3", -- 0x0F50
		x"C7",x"FF",x"FF",x"FF",x"08",x"00",x"00",x"00", -- 0x0F58
		x"FE",x"DE",x"DE",x"DF",x"C3",x"FF",x"EF",x"CF", -- 0x0F60
		x"CF",x"C0",x"C1",x"F1",x"E1",x"E3",x"FF",x"FF", -- 0x0F68
		x"0C",x"08",x"18",x"F8",x"BF",x"BB",x"BB",x"8B", -- 0x0F70
		x"98",x"FF",x"7B",x"7B",x"7B",x"09",x"FF",x"FF", -- 0x0F78
		x"FF",x"FF",x"EF",x"CF",x"CF",x"C0",x"C0",x"FF", -- 0x0F80
		x"DF",x"DF",x"C7",x"FB",x"DB",x"DB",x"D8",x"CC", -- 0x0F88
		x"FF",x"E1",x"C1",x"C1",x"C1",x"43",x"FF",x"7F", -- 0x0F90
		x"7F",x"07",x"FF",x"F7",x"F7",x"F7",x"17",x"73", -- 0x0F98
		x"E0",x"C0",x"C8",x"FF",x"EF",x"EF",x"EF",x"E0", -- 0x0FA0
		x"FF",x"EF",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF", -- 0x0FA8
		x"7F",x"3F",x"BF",x"BF",x"83",x"FF",x"DF",x"DF", -- 0x0FB0
		x"DF",x"DF",x"C3",x"E1",x"41",x"C3",x"FF",x"FF", -- 0x0FB8
		x"FF",x"FF",x"EF",x"CF",x"CF",x"CC",x"C0",x"CE", -- 0x0FC0
		x"FF",x"FF",x"E3",x"C3",x"C2",x"C6",x"FE",x"DE", -- 0x0FC8
		x"FF",x"FF",x"77",x"E7",x"E7",x"67",x"23",x"67", -- 0x0FD0
		x"FF",x"FF",x"FF",x"7F",x"7F",x"7F",x"03",x"07", -- 0x0FD8
		x"DF",x"C5",x"FD",x"FD",x"FC",x"FF",x"E7",x"C7", -- 0x0FE0
		x"C7",x"C7",x"C3",x"CB",x"FB",x"F8",x"FF",x"FF", -- 0x0FE8
		x"EF",x"EF",x"EF",x"E3",x"3F",x"DF",x"DF",x"DF", -- 0x0FF0
		x"C3",x"F9",x"F1",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x0FF8
		x"FF",x"FF",x"FF",x"DF",x"DF",x"DF",x"DF",x"C3", -- 0x1000
		x"FF",x"FF",x"FF",x"FE",x"FC",x"FC",x"FC",x"FF", -- 0x1008
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"87",x"FF", -- 0x1010
		x"FF",x"FF",x"F9",x"11",x"11",x"11",x"33",x"FF", -- 0x1018
		x"FF",x"FF",x"FF",x"DF",x"DF",x"C7",x"FF",x"FF", -- 0x1020
		x"FF",x"FF",x"FF",x"EF",x"EF",x"EF",x"E1",x"FF", -- 0x1028
		x"FF",x"FF",x"FF",x"DF",x"DF",x"DF",x"CF",x"FF", -- 0x1030
		x"FF",x"FF",x"F9",x"F1",x"F1",x"F1",x"F3",x"FF", -- 0x1038
		x"FF",x"FF",x"FF",x"DF",x"DF",x"C3",x"FF",x"FF", -- 0x1040
		x"FF",x"FF",x"DF",x"DF",x"DF",x"C7",x"FF",x"FF", -- 0x1048
		x"FF",x"EF",x"EF",x"E3",x"FF",x"FF",x"FF",x"FF", -- 0x1050
		x"FF",x"FF",x"FF",x"BF",x"BF",x"BF",x"87",x"FF", -- 0x1058
		x"FF",x"FF",x"FF",x"DF",x"DF",x"DF",x"C1",x"FF", -- 0x1060
		x"FF",x"DF",x"DF",x"DF",x"DF",x"CF",x"FF",x"FF", -- 0x1068
		x"FF",x"FF",x"FF",x"EF",x"EF",x"EF",x"E7",x"FF", -- 0x1070
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1078
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"FF", -- 0x1080
		x"9F",x"1F",x"1F",x"1F",x"2F",x"EF",x"E3",x"FF", -- 0x1088
		x"FF",x"FF",x"FF",x"7F",x"7F",x"0F",x"FF",x"FF", -- 0x1090
		x"FF",x"FF",x"FF",x"BF",x"BF",x"87",x"FF",x"FF", -- 0x1098
		x"FF",x"E7",x"C7",x"C7",x"C7",x"CF",x"FF",x"FF", -- 0x10A0
		x"FF",x"FF",x"EF",x"EF",x"EF",x"E1",x"FF",x"FF", -- 0x10A8
		x"FF",x"FF",x"FF",x"7F",x"7F",x"7F",x"03",x"FF", -- 0x10B0
		x"FF",x"FF",x"FF",x"FF",x"87",x"07",x"07",x"0F", -- 0x10B8
		x"FF",x"FF",x"FE",x"BE",x"BE",x"BF",x"9F",x"FF", -- 0x10C0
		x"FF",x"FF",x"EE",x"EE",x"EE",x"E6",x"FF",x"FF", -- 0x10C8
		x"FF",x"FF",x"FF",x"FF",x"3F",x"FF",x"FF",x"FF", -- 0x10D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"FF",x"FF", -- 0x10D8
		x"FF",x"FF",x"E3",x"C3",x"C3",x"C3",x"C7",x"FF", -- 0x10E0
		x"FF",x"FF",x"FF",x"BF",x"BF",x"87",x"FF",x"FF", -- 0x10E8
		x"FF",x"FF",x"BF",x"BF",x"8F",x"FF",x"FF",x"FF", -- 0x10F0
		x"FF",x"FF",x"FF",x"BF",x"BF",x"8F",x"FF",x"FF", -- 0x10F8
		x"FF",x"FF",x"EF",x"E1",x"FF",x"FF",x"FF",x"7F", -- 0x1100
		x"7F",x"7F",x"7F",x"0F",x"FF",x"FF",x"FF",x"FF", -- 0x1108
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"E3", -- 0x1110
		x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"07",x"FF", -- 0x1118
		x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"F8",x"FF", -- 0x1120
		x"FF",x"FF",x"FF",x"FF",x"8F",x"0F",x"0F",x"1F", -- 0x1128
		x"FF",x"FF",x"FF",x"F7",x"F7",x"F7",x"77",x"F3", -- 0x1130
		x"FF",x"FF",x"BF",x"BF",x"BF",x"87",x"FF",x"FF", -- 0x1138
		x"FF",x"FF",x"BF",x"BF",x"BF",x"BF",x"8F",x"FF", -- 0x1140
		x"FF",x"FF",x"FF",x"C7",x"87",x"8F",x"FF",x"FF", -- 0x1148
		x"FF",x"FF",x"7F",x"7F",x"0F",x"FF",x"FF",x"FF", -- 0x1150
		x"FF",x"FF",x"EF",x"EF",x"EF",x"E7",x"FF",x"FF", -- 0x1158
		x"FF",x"FF",x"FF",x"BF",x"BF",x"BF",x"BF",x"9F", -- 0x1160
		x"FF",x"FF",x"FF",x"FF",x"DF",x"DF",x"C7",x"FF", -- 0x1168
		x"FF",x"FF",x"FF",x"BF",x"BF",x"BF",x"BF",x"8F", -- 0x1170
		x"FF",x"FF",x"FF",x"DF",x"C7",x"FF",x"FF",x"FF", -- 0x1178
		x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"EF",x"EF", -- 0x1180
		x"E3",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF", -- 0x1188
		x"FF",x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF", -- 0x1190
		x"FF",x"FF",x"FF",x"FF",x"0F",x"FF",x"FF",x"FF", -- 0x1198
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x11A0
		x"FC",x"F8",x"F8",x"F8",x"FF",x"FF",x"FF",x"FF", -- 0x11A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11B0
		x"2F",x"3F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x11B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"F7",x"F7", -- 0x11C0
		x"F1",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x11C8
		x"FF",x"FF",x"FF",x"DF",x"C3",x"FF",x"FF",x"FF", -- 0x11D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11D8
		x"FF",x"FF",x"FF",x"BF",x"BF",x"87",x"FF",x"FF", -- 0x11E0
		x"FF",x"E6",x"C6",x"C6",x"C6",x"C7",x"CF",x"FF", -- 0x11E8
		x"FF",x"FF",x"FF",x"FF",x"F7",x"F7",x"F7",x"F3", -- 0x11F0
		x"FF",x"FF",x"FF",x"FF",x"3F",x"F7",x"FF",x"FF", -- 0x11F8
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FE",x"FF", -- 0x1200
		x"FF",x"FF",x"FF",x"1F",x"1F",x"9B",x"87",x"87", -- 0x1208
		x"FF",x"FF",x"3F",x"53",x"1B",x"3F",x"17",x"07", -- 0x1210
		x"87",x"8F",x"9F",x"9F",x"FF",x"FF",x"C7",x"E7", -- 0x1218
		x"82",x"89",x"8D",x"82",x"86",x"83",x"91",x"97", -- 0x1220
		x"9F",x"83",x"86",x"83",x"83",x"F3",x"FF",x"73", -- 0x1228
		x"E7",x"E7",x"E7",x"FF",x"7F",x"FF",x"C3",x"C3", -- 0x1230
		x"73",x"F3",x"F3",x"F3",x"F3",x"FF",x"FF",x"FF", -- 0x1238
		x"5C",x"3C",x"FF",x"AF",x"1F",x"7F",x"FF",x"63", -- 0x1240
		x"E3",x"F3",x"F3",x"F3",x"33",x"33",x"F3",x"FF", -- 0x1248
		x"03",x"03",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3", -- 0x1250
		x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"FF",x"FF", -- 0x1258
		x"FF",x"FF",x"FF",x"00",x"00",x"FC",x"FF",x"FD", -- 0x1260
		x"F7",x"65",x"E3",x"00",x"C1",x"E7",x"FF",x"FF", -- 0x1268
		x"FF",x"FF",x"FF",x"9F",x"9F",x"37",x"0F",x"1F", -- 0x1270
		x"8F",x"9D",x"17",x"17",x"07",x"9F",x"FF",x"FF", -- 0x1278
		x"FF",x"FF",x"7F",x"3F",x"00",x"00",x"FF",x"FF", -- 0x1280
		x"9F",x"9F",x"99",x"93",x"83",x"E1",x"E0",x"F0", -- 0x1288
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF", -- 0x1290
		x"FF",x"FB",x"E7",x"C7",x"E9",x"77",x"EE",x"5E", -- 0x1298
		x"00",x"00",x"F0",x"FC",x"9C",x"9B",x"97",x"81", -- 0x12A0
		x"EA",x"CC",x"9C",x"84",x"80",x"E6",x"00",x"00", -- 0x12A8
		x"1C",x"0E",x"57",x"6F",x"B7",x"7D",x"FD",x"DD", -- 0x12B0
		x"5D",x"ED",x"DC",x"3F",x"3F",x"1B",x"07",x"03", -- 0x12B8
		x"FF",x"BF",x"9F",x"9F",x"9E",x"92",x"93",x"90", -- 0x12C0
		x"80",x"81",x"81",x"F0",x"F0",x"B9",x"5B",x"7C", -- 0x12C8
		x"25",x"DD",x"9D",x"0C",x"3E",x"1F",x"1F",x"0F", -- 0x12D0
		x"BF",x"9B",x"FF",x"EB",x"E7",x"57",x"9B",x"91", -- 0x12D8
		x"B7",x"2F",x"07",x"0B",x"03",x"0E",x"00",x"03", -- 0x12E0
		x"FF",x"DF",x"F7",x"2F",x"03",x"07",x"83",x"E7", -- 0x12E8
		x"8B",x"08",x"81",x"C8",x"C0",x"0F",x"7F",x"FF", -- 0x12F0
		x"FF",x"F7",x"E7",x"AE",x"16",x"07",x"9F",x"FF", -- 0x12F8
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FE",x"FE", -- 0x1300
		x"FF",x"FF",x"DF",x"DF",x"EF",x"7F",x"FB",x"57", -- 0x1308
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"7F",x"7F", -- 0x1310
		x"FF",x"FF",x"FF",x"80",x"80",x"FF",x"FF",x"FF", -- 0x1318
		x"3F",x"0F",x"20",x"C0",x"5F",x"41",x"7F",x"7F", -- 0x1320
		x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"EF",x"AF", -- 0x1328
		x"FF",x"FF",x"EF",x"AF",x"AF",x"AF",x"E7",x"67", -- 0x1330
		x"67",x"67",x"67",x"67",x"67",x"0F",x"AF",x"AF", -- 0x1338
		x"A0",x"BF",x"80",x"FF",x"F5",x"EB",x"C2",x"81", -- 0x1340
		x"80",x"E7",x"E7",x"E7",x"FF",x"FF",x"D7",x"CF", -- 0x1348
		x"0D",x"FB",x"12",x"F1",x"F0",x"B3",x"83",x"A1", -- 0x1350
		x"20",x"91",x"CF",x"E7",x"F0",x"F8",x"FF",x"FF", -- 0x1358
		x"0F",x"83",x"E7",x"00",x"00",x"FF",x"FF",x"FF", -- 0x1360
		x"FF",x"FB",x"DF",x"17",x"09",x"04",x"C7",x"FF", -- 0x1368
		x"FF",x"FF",x"FF",x"00",x"00",x"F7",x"EB",x"C7", -- 0x1370
		x"CF",x"EB",x"F4",x"5B",x"20",x"01",x"11",x"FF", -- 0x1378
		x"FF",x"FF",x"FF",x"F7",x"CE",x"CB",x"D7",x"8A", -- 0x1380
		x"80",x"C6",x"C7",x"E7",x"E2",x"E1",x"E6",x"EC", -- 0x1388
		x"FF",x"FF",x"DF",x"BF",x"B6",x"5B",x"39",x"0F", -- 0x1390
		x"0F",x"1F",x"C1",x"C1",x"FF",x"FF",x"E7",x"E7", -- 0x1398
		x"C7",x"E7",x"E3",x"F3",x"FF",x"FF",x"F0",x"F0", -- 0x13A0
		x"FF",x"FF",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC", -- 0x13A8
		x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F", -- 0x13B0
		x"CF",x"FF",x"FF",x"CF",x"DF",x"3F",x"2F",x"5F", -- 0x13B8
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC", -- 0x13C0
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC", -- 0x13C8
		x"15",x"2F",x"3F",x"1B",x"17",x"07",x"8F",x"9F", -- 0x13D0
		x"E1",x"E0",x"FF",x"FF",x"FB",x"F3",x"F3",x"F3", -- 0x13D8
		x"F7",x"E7",x"E3",x"F5",x"EB",x"E7",x"C6",x"C9", -- 0x13E0
		x"CA",x"C1",x"E5",x"E0",x"F0",x"FB",x"FF",x"FF", -- 0x13E8
		x"F0",x"F0",x"F0",x"F2",x"F2",x"F3",x"F0",x"F0", -- 0x13F0
		x"FF",x"FE",x"7C",x"2F",x"15",x"03",x"C3",x"FF", -- 0x13F8
		x"55",x"A4",x"A9",x"44",x"53",x"A9",x"15",x"FF", -- 0x1400
		x"6B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1408
		x"55",x"CB",x"AD",x"CB",x"AA",x"77",x"21",x"CA", -- 0x1410
		x"BF",x"AD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1418
		x"B4",x"15",x"A4",x"8B",x"36",x"96",x"CD",x"4C", -- 0x1420
		x"15",x"EA",x"3F",x"2B",x"80",x"FF",x"FF",x"FF", -- 0x1428
		x"55",x"44",x"A9",x"6B",x"D0",x"6B",x"45",x"AA", -- 0x1430
		x"52",x"A2",x"D5",x"FF",x"1E",x"80",x"FF",x"FF", -- 0x1438
		x"C0",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1440
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1448
		x"03",x"03",x"03",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1450
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1458
		x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1460
		x"FF",x"FF",x"FF",x"FF",x"FD",x"F9",x"F9",x"FB", -- 0x1468
		x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1470
		x"FF",x"FF",x"FF",x"FF",x"FF",x"E3",x"CF",x"57", -- 0x1478
		x"B5",x"4A",x"3A",x"AD",x"0B",x"51",x"C4",x"3E", -- 0x1480
		x"43",x"B8",x"4C",x"A8",x"CA",x"8E",x"E6",x"EB", -- 0x1488
		x"55",x"6A",x"B0",x"9D",x"49",x"36",x"91",x"3D", -- 0x1490
		x"46",x"39",x"75",x"C5",x"B9",x"CD",x"EC",x"7C", -- 0x1498
		x"00",x"01",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14A8
		x"00",x"55",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14B8
		x"AA",x"A5",x"94",x"56",x"34",x"C9",x"EE",x"D3", -- 0x14C0
		x"75",x"7D",x"BB",x"DC",x"EC",x"F7",x"F7",x"FB", -- 0x14C8
		x"AA",x"71",x"1A",x"DD",x"29",x"D2",x"FC",x"2B", -- 0x14D0
		x"55",x"6E",x"15",x"79",x"CE",x"4D",x"54",x"25", -- 0x14D8
		x"FD",x"FE",x"FE",x"FF",x"FF",x"FF",x"0F",x"3F", -- 0x14E0
		x"3F",x"0F",x"FF",x"83",x"9B",x"9B",x"9B",x"9B", -- 0x14E8
		x"AE",x"F5",x"D6",x"6F",x"7B",x"B4",x"FA",x"DB", -- 0x14F0
		x"EF",x"EC",x"EF",x"F7",x"F6",x"FB",x"FB",x"FB", -- 0x14F8
		x"AA",x"6C",x"93",x"6A",x"D0",x"26",x"55",x"FF", -- 0x1500
		x"AA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1508
		x"AA",x"55",x"52",x"F4",x"AF",x"A5",x"2D",x"FF", -- 0x1510
		x"DD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1518
		x"AA",x"55",x"D5",x"AB",x"65",x"94",x"CA",x"52", -- 0x1520
		x"5B",x"FF",x"AE",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1528
		x"AA",x"44",x"F5",x"A9",x"5A",x"56",x"85",x"69", -- 0x1530
		x"55",x"FF",x"BA",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1538
		x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1540
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1548
		x"F8",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8", -- 0x1550
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x1558
		x"55",x"AB",x"AE",x"57",x"00",x"55",x"FF",x"FF", -- 0x1560
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1568
		x"4B",x"55",x"B6",x"AB",x"3C",x"00",x"D5",x"FF", -- 0x1570
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1578
		x"AA",x"62",x"98",x"4F",x"B9",x"56",x"D5",x"3A", -- 0x1580
		x"D9",x"44",x"32",x"99",x"C5",x"19",x"4D",x"D1", -- 0x1588
		x"AA",x"D5",x"A9",x"B2",x"16",x"E9",x"DC",x"35", -- 0x1590
		x"58",x"7F",x"C1",x"BD",x"D5",x"7D",x"D5",x"E5", -- 0x1598
		x"FE",x"00",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15A8
		x"00",x"00",x"AA",x"FF",x"F8",x"F8",x"F8",x"F8", -- 0x15B0
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x15B8
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15C8
		x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x15D0
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x15D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E8
		x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD", -- 0x15F0
		x"BD",x"BF",x"BF",x"BF",x"BF",x"FF",x"FF",x"FF", -- 0x15F8
		x"AA",x"55",x"26",x"2A",x"00",x"FF",x"41",x"FF", -- 0x1600
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1608
		x"AB",x"44",x"56",x"A9",x"25",x"EE",x"3F",x"84", -- 0x1610
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1618
		x"AA",x"14",x"B5",x"D2",x"67",x"59",x"AA",x"55", -- 0x1620
		x"D5",x"7F",x"15",x"C0",x"FF",x"FF",x"FF",x"FF", -- 0x1628
		x"AA",x"55",x"35",x"C4",x"2B",x"B6",x"49",x"5B", -- 0x1630
		x"54",x"FF",x"6B",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1640
		x"FF",x"FE",x"FC",x"F8",x"E0",x"C2",x"05",x"0A", -- 0x1648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"F8",x"F0", -- 0x1650
		x"81",x"02",x"09",x"36",x"C8",x"17",x"29",x"A6", -- 0x1658
		x"66",x"84",x"01",x"C4",x"EE",x"FF",x"FF",x"FF", -- 0x1660
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1668
		x"EB",x"E5",x"0A",x"63",x"F0",x"E5",x"FF",x"F8", -- 0x1670
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x1678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1680
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1688
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1690
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1698
		x"AA",x"5D",x"00",x"AA",x"FF",x"FF",x"FF",x"FF", -- 0x16A0
		x"FF",x"FF",x"FF",x"FF",x"FD",x"F9",x"F9",x"FB", -- 0x16A8
		x"00",x"00",x"2A",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"E3",x"CF",x"57", -- 0x16B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16C8
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x16D0
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x16D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16E8
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x16F0
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x16F8
		x"AA",x"54",x"E5",x"99",x"80",x"3F",x"4E",x"9F", -- 0x1700
		x"7F",x"5F",x"7F",x"5F",x"7F",x"5F",x"7F",x"5F", -- 0x1708
		x"AA",x"B5",x"6C",x"C9",x"00",x"FF",x"BA",x"FF", -- 0x1710
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1718
		x"BA",x"4B",x"35",x"4A",x"A8",x"91",x"A4",x"5B", -- 0x1720
		x"FF",x"BA",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1728
		x"AA",x"55",x"34",x"9A",x"A5",x"56",x"55",x"6D", -- 0x1730
		x"FF",x"EB",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1738
		x"AA",x"13",x"B5",x"2A",x"B6",x"D5",x"DD",x"45", -- 0x1740
		x"AA",x"00",x"75",x"FF",x"51",x"00",x"FE",x"FF", -- 0x1748
		x"AA",x"11",x"6E",x"9D",x"A3",x"56",x"2B",x"EA", -- 0x1750
		x"93",x"5D",x"32",x"A9",x"FC",x"E6",x"00",x"FE", -- 0x1758
		x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1760
		x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"9E",x"8C", -- 0x1768
		x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x1778
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1788
		x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1790
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1798
		x"AA",x"54",x"9A",x"24",x"01",x"57",x"FF",x"FF", -- 0x17A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"9E",x"8C", -- 0x17A8
		x"AA",x"D5",x"44",x"00",x"55",x"FF",x"FF",x"FF", -- 0x17B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x17B8
		x"B5",x"6A",x"5F",x"9B",x"BE",x"2A",x"55",x"D4", -- 0x17C0
		x"21",x"D7",x"1F",x"3F",x"7F",x"FF",x"FF",x"FF", -- 0x17C8
		x"75",x"AA",x"DA",x"74",x"A6",x"D4",x"24",x"98", -- 0x17D0
		x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x17D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E8
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x17F0
		x"F8",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1800
		x"FF",x"FF",x"FF",x"00",x"AA",x"00",x"FF",x"FF", -- 0x1808
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1810
		x"FF",x"FF",x"FF",x"7F",x"80",x"2A",x"80",x"BD", -- 0x1818
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1820
		x"FF",x"00",x"56",x"01",x"FC",x"FF",x"FF",x"FF", -- 0x1828
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1830
		x"FF",x"FF",x"00",x"55",x"00",x"FF",x"FF",x"FF", -- 0x1838
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1840
		x"FF",x"00",x"55",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1848
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1850
		x"00",x"55",x"00",x"3F",x"FF",x"FF",x"FF",x"FF", -- 0x1858
		x"7F",x"5F",x"7F",x"5F",x"7F",x"5F",x"7F",x"1F", -- 0x1860
		x"00",x"3B",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1868
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1870
		x"00",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1878
		x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"DF",x"EF", -- 0x1880
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"03", -- 0x1888
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x1890
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x1898
		x"7F",x"3F",x"47",x"3F",x"3F",x"1F",x"0F",x"0F", -- 0x18A0
		x"0F",x"0F",x"3F",x"08",x"CE",x"C9",x"9C",x"FF", -- 0x18A8
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x18B0
		x"F8",x"FF",x"C5",x"E0",x"73",x"0B",x"E7",x"FF", -- 0x18B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
		x"01",x"FD",x"BD",x"7D",x"7D",x"35",x"8D",x"7F", -- 0x18E0
		x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E8
		x"01",x"FD",x"DD",x"5D",x"5D",x"65",x"7D",x"1E", -- 0x18F0
		x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F8
		x"55",x"AB",x"AE",x"57",x"D5",x"2B",x"53",x"D5", -- 0x1900
		x"2B",x"55",x"03",x"54",x"FD",x"FF",x"FF",x"FF", -- 0x1908
		x"4B",x"55",x"B6",x"AB",x"7C",x"77",x"BB",x"AA", -- 0x1910
		x"65",x"7D",x"DE",x"0A",x"50",x"F5",x"FF",x"F8", -- 0x1918
		x"FF",x"FF",x"FF",x"07",x"03",x"01",x"00",x"00", -- 0x1920
		x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0", -- 0x1928
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"78", -- 0x1930
		x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"38", -- 0x1938
		x"20",x"20",x"20",x"E0",x"C0",x"80",x"00",x"00", -- 0x1940
		x"00",x"00",x"01",x"03",x"07",x"FF",x"FF",x"FF", -- 0x1948
		x"28",x"28",x"28",x"38",x"38",x"38",x"38",x"38", -- 0x1950
		x"78",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x1958
		x"FF",x"FF",x"F8",x"01",x"54",x"03",x"C3",x"C6", -- 0x1960
		x"86",x"8D",x"0B",x"16",x"1D",x"36",x"1A",x"EB", -- 0x1968
		x"F8",x"E0",x"05",x"50",x"0C",x"7B",x"4D",x"B2", -- 0x1970
		x"97",x"B5",x"6A",x"AD",x"AB",x"D6",x"B5",x"4B", -- 0x1978
		x"FF",x"FF",x"FF",x"83",x"18",x"18",x"9F",x"FF", -- 0x1980
		x"0F",x"EE",x"EC",x"E9",x"70",x"70",x"30",x"B0", -- 0x1988
		x"FF",x"FF",x"FF",x"C1",x"8D",x"0E",x"CF",x"FF", -- 0x1990
		x"FF",x"E3",x"F9",x"FD",x"01",x"01",x"08",x"C0", -- 0x1998
		x"F0",x"F1",x"F0",x"30",x"30",x"38",x"7C",x"EE", -- 0x19A0
		x"CF",x"98",x"32",x"70",x"60",x"00",x"00",x"00", -- 0x19A8
		x"01",x"FE",x"7E",x"1D",x"01",x"03",x"05",x"FC", -- 0x19B0
		x"F0",x"E0",x"C0",x"00",x"01",x"01",x"01",x"01", -- 0x19B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D8
		x"01",x"03",x"03",x"02",x"02",x"03",x"01",x"00", -- 0x19E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E8
		x"01",x"55",x"55",x"95",x"D1",x"49",x"9F",x"FE", -- 0x19F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F8
		x"55",x"AB",x"AE",x"57",x"D5",x"2B",x"D5",x"00", -- 0x1A00
		x"80",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A08
		x"4B",x"55",x"B6",x"AB",x"7C",x"77",x"BB",x"AA", -- 0x1A10
		x"00",x"00",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A18
		x"FF",x"FF",x"FF",x"0F",x"07",x"03",x"00",x"00", -- 0x1A20
		x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0", -- 0x1A28
		x"FF",x"FF",x"FF",x"C0",x"80",x"00",x"00",x"00", -- 0x1A30
		x"00",x"00",x"07",x"0F",x"1F",x"1F",x"1F",x"1F", -- 0x1A38
		x"20",x"20",x"20",x"E0",x"C0",x"80",x"00",x"00", -- 0x1A40
		x"00",x"00",x"03",x"07",x"0F",x"FF",x"FF",x"FF", -- 0x1A48
		x"10",x"10",x"10",x"1F",x"0F",x"07",x"00",x"00", -- 0x1A50
		x"00",x"00",x"00",x"80",x"C0",x"FF",x"FF",x"FF", -- 0x1A58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"2A",x"80", -- 0x1A60
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A68
		x"FF",x"FF",x"FF",x"FF",x"80",x"2A",x"00",x"FF", -- 0x1A70
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F0",x"E0", -- 0x1A78
		x"97",x"18",x"FC",x"FF",x"FF",x"00",x"FF",x"FF", -- 0x1A80
		x"BB",x"BF",x"07",x"31",x"03",x"07",x"06",x"06", -- 0x1A88
		x"FF",x"FF",x"7F",x"7F",x"7F",x"FF",x"FF",x"FF", -- 0x1A90
		x"FC",x"FF",x"FF",x"E1",x"FC",x"FF",x"83",x"73", -- 0x1A98
		x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA0
		x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AA8
		x"2B",x"1B",x"0F",x"07",x"03",x"06",x"00",x"00", -- 0x1AB0
		x"01",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD8
		x"F9",x"F3",x"F1",x"F4",x"FE",x"FC",x"FC",x"F9", -- 0x1AE0
		x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AE8
		x"FF",x"C7",x"9F",x"AF",x"1F",x"4F",x"BF",x"5F", -- 0x1AF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AF8
		x"55",x"AB",x"AE",x"57",x"D5",x"04",x"50",x"F5", -- 0x1B00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B08
		x"4B",x"55",x"B6",x"AB",x"7C",x"AA",x"34",x"00", -- 0x1B10
		x"D5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8", -- 0x1B20
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x1B28
		x"FF",x"FF",x"FF",x"80",x"00",x"00",x"00",x"00", -- 0x1B30
		x"00",x"00",x"07",x"0F",x"1F",x"1F",x"1F",x"1F", -- 0x1B38
		x"10",x"10",x"10",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x1B40
		x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B48
		x"10",x"10",x"10",x"1F",x"0F",x"07",x"00",x"00", -- 0x1B50
		x"00",x"00",x"00",x"00",x"80",x"FF",x"FF",x"FF", -- 0x1B58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0", -- 0x1B60
		x"05",x"50",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"55", -- 0x1B70
		x"00",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B78
		x"FF",x"00",x"FF",x"FF",x"7F",x"1E",x"06",x"C0", -- 0x1B80
		x"3C",x"06",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x1B88
		x"FF",x"00",x"FF",x"00",x"E4",x"C6",x"C6",x"C7", -- 0x1B90
		x"C0",x"40",x"80",x"9C",x"DE",x"4F",x"41",x"41", -- 0x1B98
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"0C", -- 0x1BA0
		x"F0",x"01",x"03",x"E1",x"00",x"00",x"00",x"00", -- 0x1BA8
		x"41",x"41",x"41",x"81",x"83",x"03",x"03",x"02", -- 0x1BB0
		x"00",x"80",x"C0",x"C0",x"8C",x"00",x"00",x"00", -- 0x1BB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BE0
		x"1F",x"0F",x"03",x"00",x"00",x"A0",x"D0",x"54", -- 0x1BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF0
		x"FF",x"FF",x"FF",x"3F",x"1F",x"0F",x"01",x"00", -- 0x1BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x1FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
