-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_A6 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_A6 is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"20",x"48",x"50",x"71",x"77",x"A9",x"72",x"39", -- 0x0000
		x"7B",x"7E",x"AC",x"5D",x"6E",x"3A",x"31",x"21", -- 0x0008
		x"FF",x"7F",x"BF",x"4F",x"83",x"03",x"83",x"09", -- 0x0010
		x"8C",x"D1",x"F2",x"DF",x"6E",x"F9",x"56",x"30", -- 0x0018
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0020
		x"7F",x"1F",x"47",x"C7",x"43",x"E9",x"79",x"A0", -- 0x0028
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0030
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0038
		x"10",x"B0",x"64",x"2A",x"4E",x"B4",x"FC",x"70", -- 0x0040
		x"15",x"AA",x"22",x"C5",x"F6",x"6E",x"3D",x"91", -- 0x0048
		x"7F",x"7F",x"7F",x"7F",x"FF",x"7F",x"3F",x"1F", -- 0x0050
		x"1F",x"0F",x"07",x"87",x"B7",x"6F",x"DF",x"1F", -- 0x0058
		x"00",x"20",x"F2",x"AB",x"76",x"9F",x"81",x"E0", -- 0x0060
		x"D5",x"7B",x"BC",x"5A",x"0C",x"12",x"21",x"19", -- 0x0068
		x"BF",x"DF",x"3F",x"7F",x"3F",x"1F",x"9F",x"1F", -- 0x0070
		x"BF",x"3F",x"7F",x"7F",x"3F",x"3F",x"1F",x"1F", -- 0x0078
		x"4C",x"B9",x"FA",x"EF",x"27",x"83",x"99",x"D0", -- 0x0080
		x"7A",x"3C",x"F9",x"93",x"B3",x"E7",x"EF",x"CF", -- 0x0088
		x"1F",x"1F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0090
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0098
		x"DF",x"9F",x"1F",x"0F",x"4F",x"8F",x"5F",x"9F", -- 0x00A0
		x"3F",x"3F",x"1F",x"9F",x"8F",x"CF",x"EF",x"4F", -- 0x00A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B8
		x"0F",x"8F",x"87",x"C7",x"27",x"CF",x"8F",x"1F", -- 0x00C0
		x"0F",x"47",x"83",x"DB",x"F1",x"E1",x"40",x"10", -- 0x00C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D8
		x"10",x"A8",x"F1",x"F1",x"28",x"50",x"CC",x"00", -- 0x00E0
		x"B4",x"59",x"0B",x"DF",x"B5",x"F1",x"78",x"10", -- 0x00E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F", -- 0x00F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F8
		x"10",x"B8",x"E9",x"A9",x"03",x"87",x"CF",x"CF", -- 0x0100
		x"A7",x"47",x"83",x"83",x"A3",x"53",x"07",x"CF", -- 0x0108
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0110
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0118
		x"20",x"51",x"AE",x"DC",x"7E",x"E9",x"50",x"0A", -- 0x0120
		x"1B",x"5D",x"AF",x"47",x"63",x"62",x"F0",x"92", -- 0x0128
		x"0F",x"0F",x"9F",x"3F",x"3F",x"9F",x"8F",x"0F", -- 0x0130
		x"6F",x"0F",x"DF",x"9F",x"FF",x"7F",x"FF",x"FF", -- 0x0138
		x"02",x"C8",x"B5",x"C9",x"B9",x"E3",x"CF",x"3F", -- 0x0140
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0148
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0150
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0158
		x"00",x"22",x"22",x"56",x"6F",x"15",x"9C",x"FE", -- 0x0160
		x"77",x"0A",x"2C",x"36",x"BC",x"5F",x"67",x"00", -- 0x0168
		x"FF",x"7F",x"3F",x"3F",x"3C",x"38",x"00",x"82", -- 0x0170
		x"B4",x"5C",x"72",x"E8",x"38",x"F2",x"3E",x"0C", -- 0x0178
		x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"1F", -- 0x0180
		x"0F",x"0F",x"9F",x"8F",x"83",x"61",x"50",x"B0", -- 0x0188
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0190
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0198
		x"10",x"B8",x"EE",x"ED",x"34",x"80",x"80",x"44", -- 0x01A0
		x"23",x"CF",x"9F",x"3F",x"FF",x"FF",x"FF",x"FF", -- 0x01A8
		x"0F",x"8F",x"3F",x"FF",x"FF",x"7F",x"7F",x"FF", -- 0x01B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01B8
		x"C0",x"20",x"93",x"0C",x"05",x"52",x"44",x"2C", -- 0x01C0
		x"20",x"1A",x"0E",x"B3",x"0D",x"15",x"88",x"42", -- 0x01C8
		x"08",x"54",x"24",x"9A",x"AD",x"FA",x"51",x"24", -- 0x01D0
		x"1D",x"B9",x"FB",x"E3",x"83",x"17",x"7F",x"FF", -- 0x01D8
		x"FF",x"FF",x"FF",x"CF",x"83",x"20",x"A0",x"91", -- 0x01E0
		x"51",x"07",x"92",x"E1",x"B1",x"E8",x"7E",x"1C", -- 0x01E8
		x"FF",x"FF",x"FF",x"F9",x"E0",x"D0",x"30",x"39", -- 0x01F0
		x"B4",x"AA",x"1D",x"04",x"98",x"E6",x"EB",x"00", -- 0x01F8
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"9C",x"02", -- 0x0200
		x"64",x"46",x"A3",x"A1",x"93",x"69",x"54",x"B0", -- 0x0208
		x"FF",x"FF",x"F1",x"C1",x"00",x"20",x"28",x"32", -- 0x0210
		x"51",x"82",x"48",x"40",x"64",x"F9",x"56",x"30", -- 0x0218
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0220
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0228
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0230
		x"FC",x"F1",x"C2",x"C5",x"92",x"A0",x"36",x"64", -- 0x0238
		x"FF",x"FF",x"FC",x"F8",x"FA",x"F2",x"F4",x"F7", -- 0x0240
		x"F3",x"FB",x"F8",x"F0",x"F0",x"F0",x"F3",x"F4", -- 0x0248
		x"36",x"6C",x"2A",x"1E",x"1D",x"8C",x"A2",x"54", -- 0x0250
		x"80",x"C8",x"C8",x"64",x"95",x"4A",x"A0",x"D8", -- 0x0258
		x"F7",x"F5",x"E4",x"CE",x"D8",x"B5",x"9A",x"B3", -- 0x0260
		x"A8",x"B8",x"D6",x"D4",x"E8",x"ED",x"F2",x"F6", -- 0x0268
		x"A0",x"18",x"54",x"40",x"20",x"42",x"E8",x"94", -- 0x0270
		x"00",x"48",x"C8",x"64",x"95",x"8A",x"20",x"D8", -- 0x0278
		x"E7",x"F6",x"F2",x"FB",x"F9",x"FD",x"FD",x"FC", -- 0x0280
		x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0288
		x"20",x"18",x"94",x"D8",x"00",x"82",x"A8",x"D4", -- 0x0290
		x"B8",x"7C",x"68",x"A4",x"95",x"AA",x"20",x"58", -- 0x0298
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02A8
		x"26",x"AC",x"8A",x"CE",x"CD",x"E4",x"F9",x"FE", -- 0x02B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02B8
		x"00",x"A1",x"E8",x"69",x"37",x"88",x"E0",x"39", -- 0x02C0
		x"D1",x"F8",x"EC",x"F7",x"F1",x"FD",x"FE",x"FF", -- 0x02C8
		x"A0",x"98",x"D4",x"C0",x"A0",x"C2",x"28",x"14", -- 0x02D0
		x"00",x"88",x"88",x"24",x"95",x"AA",x"A0",x"58", -- 0x02D8
		x"11",x"B8",x"E8",x"EE",x"24",x"FD",x"8B",x"2E", -- 0x02E0
		x"F3",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02E8
		x"E6",x"C1",x"D0",x"1A",x"BC",x"1B",x"61",x"1C", -- 0x02F0
		x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02F8
		x"FF",x"FF",x"FF",x"FF",x"3F",x"0E",x"42",x"87", -- 0x0300
		x"62",x"8B",x"10",x"C9",x"8F",x"D6",x"40",x"10", -- 0x0308
		x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"0F",x"0F", -- 0x0310
		x"84",x"00",x"51",x"30",x"38",x"96",x"CB",x"00", -- 0x0318
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x0320
		x"70",x"01",x"90",x"D8",x"8D",x"C4",x"60",x"30", -- 0x0328
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"07", -- 0x0330
		x"04",x"20",x"19",x"04",x"58",x"B6",x"EB",x"00", -- 0x0338
		x"11",x"B8",x"EA",x"A9",x"16",x"93",x"9A",x"0C", -- 0x0340
		x"E6",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0348
		x"68",x"F4",x"E4",x"7A",x"1D",x"26",x"30",x"0E", -- 0x0350
		x"05",x"72",x"F9",x"FC",x"FF",x"FF",x"FF",x"FF", -- 0x0358
		x"10",x"AD",x"E6",x"3C",x"9A",x"CC",x"E0",x"FF", -- 0x0360
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0368
		x"16",x"39",x"10",x"1C",x"9A",x"2F",x"71",x"FC", -- 0x0370
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0378
		x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FD",x"FC", -- 0x0380
		x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE", -- 0x0388
		x"60",x"D8",x"54",x"60",x"68",x"D2",x"E8",x"94", -- 0x0390
		x"44",x"E8",x"4A",x"64",x"15",x"CA",x"E0",x"58", -- 0x0398
		x"FF",x"F8",x"F0",x"E0",x"E0",x"C0",x"80",x"80", -- 0x03A0
		x"80",x"C0",x"C0",x"E0",x"E2",x"F7",x"FF",x"FF", -- 0x03A8
		x"FF",x"7F",x"3F",x"1F",x"07",x"03",x"03",x"03", -- 0x03B0
		x"07",x"07",x"0F",x"3F",x"7F",x"FF",x"FF",x"FF", -- 0x03B8
		x"FF",x"FF",x"FF",x"FF",x"FD",x"F8",x"F8",x"F0", -- 0x03C0
		x"F0",x"F8",x"F8",x"FC",x"FF",x"FF",x"FF",x"FF", -- 0x03C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"3F", -- 0x03D0
		x"1F",x"1F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03D8
		x"FF",x"FF",x"FF",x"FC",x"F8",x"F8",x"F0",x"F0", -- 0x03E0
		x"F8",x"F8",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03E8
		x"FF",x"FF",x"3F",x"1F",x"0F",x"0F",x"07",x"07", -- 0x03F0
		x"07",x"07",x"4F",x"3F",x"FF",x"FF",x"FF",x"FF", -- 0x03F8
		x"DF",x"FF",x"F7",x"FF",x"FB",x"FF",x"FF",x"EF", -- 0x0400
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FE",x"7F", -- 0x0408
		x"34",x"AA",x"8D",x"F5",x"CB",x"E2",x"FA",x"FE", -- 0x0410
		x"FF",x"DF",x"BF",x"EF",x"FF",x"7F",x"BB",x"FF", -- 0x0418
		x"8A",x"E4",x"F5",x"FA",x"D4",x"FD",x"FE",x"EE", -- 0x0420
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FE",x"7F", -- 0x0428
		x"B4",x"AE",x"4D",x"55",x"A3",x"AA",x"44",x"56", -- 0x0430
		x"13",x"9F",x"FF",x"FF",x"FF",x"7F",x"BB",x"FF", -- 0x0438
		x"AA",x"54",x"41",x"28",x"CA",x"E4",x"F8",x"FE", -- 0x0440
		x"FE",x"FF",x"FF",x"FF",x"DB",x"FF",x"FE",x"7F", -- 0x0448
		x"B4",x"AA",x"49",x"54",x"83",x"88",x"44",x"54", -- 0x0450
		x"87",x"1F",x"FF",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x0458
		x"AA",x"54",x"55",x"BA",x"3A",x"D5",x"AD",x"2A", -- 0x0460
		x"CC",x"F9",x"FF",x"FF",x"FF",x"FF",x"FE",x"7F", -- 0x0468
		x"B4",x"AA",x"49",x"55",x"A3",x"AA",x"44",x"44", -- 0x0470
		x"9B",x"4F",x"FF",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x0478
		x"AA",x"54",x"51",x"B8",x"2A",x"D4",x"AC",x"2A", -- 0x0480
		x"D4",x"AA",x"68",x"13",x"D4",x"F3",x"FF",x"7F", -- 0x0488
		x"B4",x"AE",x"4D",x"54",x"83",x"88",x"44",x"54", -- 0x0490
		x"97",x"8F",x"1F",x"7F",x"FF",x"FF",x"FB",x"FF", -- 0x0498
		x"AA",x"54",x"55",x"AA",x"B2",x"55",x"AD",x"2A", -- 0x04A0
		x"D4",x"AA",x"2B",x"51",x"29",x"CF",x"7F",x"FF", -- 0x04A8
		x"B4",x"AE",x"4D",x"55",x"A1",x"AA",x"44",x"54", -- 0x04B0
		x"BB",x"AF",x"5F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x04B8
		x"AA",x"54",x"51",x"A0",x"1A",x"D4",x"AC",x"2A", -- 0x04C0
		x"D4",x"AA",x"48",x"52",x"2B",x"97",x"DF",x"0F", -- 0x04C8
		x"B4",x"AA",x"49",x"50",x"83",x"88",x"44",x"54", -- 0x04D0
		x"93",x"CF",x"BF",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x04D8
		x"AA",x"54",x"45",x"AA",x"2A",x"D5",x"AD",x"2A", -- 0x04E0
		x"D4",x"AA",x"4A",x"33",x"6D",x"94",x"D3",x"2A", -- 0x04E8
		x"B4",x"AE",x"4D",x"55",x"A3",x"AA",x"44",x"44", -- 0x04F0
		x"93",x"AF",x"1F",x"3F",x"7F",x"7F",x"FB",x"FF", -- 0x04F8
		x"AA",x"54",x"45",x"38",x"CA",x"F8",x"FC",x"FF", -- 0x0500
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FE",x"7F", -- 0x0508
		x"B4",x"AE",x"49",x"04",x"83",x"9F",x"7F",x"FF", -- 0x0510
		x"FF",x"FF",x"FF",x"EF",x"FF",x"7F",x"BB",x"FF", -- 0x0518
		x"AA",x"54",x"55",x"BA",x"2A",x"C5",x"AD",x"2A", -- 0x0520
		x"D4",x"AA",x"4B",x"31",x"CC",x"F1",x"FF",x"7F", -- 0x0528
		x"B4",x"AA",x"4D",x"54",x"A7",x"A7",x"4F",x"5F", -- 0x0530
		x"9F",x"BF",x"FF",x"7F",x"FF",x"FF",x"FB",x"FF", -- 0x0538
		x"AA",x"44",x"55",x"AA",x"3A",x"D5",x"AD",x"28", -- 0x0540
		x"D4",x"A9",x"67",x"5F",x"3F",x"BF",x"7E",x"FF", -- 0x0548
		x"B4",x"AE",x"4B",x"50",x"A3",x"B7",x"5F",x"3F", -- 0x0550
		x"7F",x"FF",x"FF",x"EF",x"FF",x"7F",x"BB",x"FF", -- 0x0558
		x"8A",x"E4",x"FB",x"FE",x"DF",x"FF",x"FF",x"EF", -- 0x0560
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FE",x"7F", -- 0x0568
		x"B4",x"A2",x"49",x"54",x"03",x"08",x"84",x"95", -- 0x0570
		x"DA",x"C2",x"E5",x"E4",x"F3",x"7F",x"BF",x"FF", -- 0x0578
		x"AA",x"54",x"51",x"A8",x"2A",x"D4",x"AC",x"2A", -- 0x0580
		x"D4",x"AA",x"68",x"33",x"CD",x"F9",x"FF",x"7F", -- 0x0588
		x"B4",x"AE",x"4D",x"54",x"83",x"88",x"44",x"55", -- 0x0590
		x"9A",x"82",x"21",x"54",x"63",x"1F",x"FF",x"FF", -- 0x0598
		x"DF",x"FF",x"F7",x"FF",x"DB",x"FF",x"FF",x"EF", -- 0x05A0
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FF",x"7F", -- 0x05A8
		x"F4",x"F2",x"E5",x"E5",x"FB",x"CA",x"D4",x"C5", -- 0x05B0
		x"FA",x"CA",x"E5",x"C5",x"E6",x"F3",x"F3",x"F1", -- 0x05B8
		x"DF",x"FF",x"FE",x"FE",x"DF",x"FC",x"FC",x"FE", -- 0x05C0
		x"FC",x"FC",x"FE",x"FE",x"DE",x"FE",x"FF",x"7F", -- 0x05C8
		x"34",x"2E",x"4D",x"54",x"83",x"8A",x"44",x"55", -- 0x05D0
		x"9A",x"A2",x"01",x"35",x"26",x"CB",x"2B",x"55", -- 0x05D8
		x"FA",x"F4",x"E5",x"EA",x"EA",x"D5",x"CD",x"CA", -- 0x05E0
		x"D4",x"CA",x"C9",x"E2",x"ED",x"EA",x"F6",x"73", -- 0x05E8
		x"B4",x"AA",x"49",x"55",x"A3",x"AA",x"44",x"55", -- 0x05F0
		x"9A",x"8A",x"25",x"55",x"62",x"A9",x"AB",x"55", -- 0x05F8
		x"DF",x"FF",x"F7",x"FF",x"DB",x"FF",x"FF",x"EF", -- 0x0600
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FE",x"7F", -- 0x0608
		x"F4",x"F6",x"ED",x"E4",x"E3",x"C8",x"D4",x"E5", -- 0x0610
		x"F2",x"FE",x"F9",x"FD",x"FC",x"7E",x"BE",x"FF", -- 0x0618
		x"DF",x"FF",x"FE",x"FE",x"FE",x"FD",x"FD",x"FE", -- 0x0620
		x"FC",x"FF",x"FF",x"FF",x"DB",x"FF",x"FE",x"7F", -- 0x0628
		x"34",x"2E",x"4D",x"55",x"A3",x"AA",x"44",x"55", -- 0x0630
		x"9A",x"AA",x"E5",x"F9",x"FC",x"7F",x"BE",x"FF", -- 0x0638
		x"F2",x"F4",x"E9",x"E0",x"F2",x"F4",x"F8",x"FC", -- 0x0640
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FE",x"7F", -- 0x0648
		x"B4",x"AA",x"49",x"54",x"A3",x"A8",x"44",x"55", -- 0x0650
		x"5A",x"C6",x"F1",x"F9",x"FC",x"7E",x"BE",x"FF", -- 0x0658
		x"AA",x"D4",x"E5",x"EA",x"F2",x"F5",x"FD",x"FA", -- 0x0660
		x"FF",x"FC",x"FE",x"FF",x"DF",x"FF",x"FE",x"7F", -- 0x0668
		x"B4",x"AE",x"4D",x"55",x"AB",x"AA",x"44",x"55", -- 0x0670
		x"9A",x"8A",x"25",x"B5",x"E6",x"FD",x"FE",x"FF", -- 0x0678
		x"AA",x"55",x"51",x"A8",x"2A",x"D5",x"AC",x"2A", -- 0x0680
		x"D4",x"8E",x"2A",x"50",x"4B",x"A7",x"CF",x"0F", -- 0x0688
		x"B5",x"AB",x"47",x"57",x"9F",x"0F",x"4F",x"5F", -- 0x0690
		x"BF",x"5F",x"3F",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x0698
		x"F2",x"F4",x"E5",x"EA",x"CA",x"ED",x"F9",x"FC", -- 0x06A0
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FF",x"7F", -- 0x06A8
		x"B4",x"AA",x"45",x"55",x"A3",x"AA",x"44",x"55", -- 0x06B0
		x"1A",x"8A",x"C5",x"D5",x"E6",x"E9",x"F7",x"F1", -- 0x06B8
		x"DF",x"FF",x"FE",x"FE",x"FD",x"FD",x"FD",x"FE", -- 0x06C0
		x"FF",x"FF",x"FF",x"FF",x"DB",x"FF",x"FF",x"7F", -- 0x06C8
		x"34",x"2E",x"4D",x"54",x"A3",x"A8",x"44",x"55", -- 0x06D0
		x"1A",x"82",x"E1",x"D5",x"E6",x"EB",x"FB",x"F5", -- 0x06D8
		x"DF",x"FF",x"FE",x"FE",x"DF",x"FE",x"FD",x"F9", -- 0x06E0
		x"F0",x"EA",x"C9",x"D3",x"E5",x"E6",x"F2",x"73", -- 0x06E8
		x"34",x"2E",x"4D",x"55",x"AB",x"AA",x"44",x"55", -- 0x06F0
		x"9A",x"8A",x"25",x"55",x"22",x"A9",x"EB",x"55", -- 0x06F8
		x"AA",x"54",x"51",x"A8",x"2A",x"D4",x"AC",x"2A", -- 0x0700
		x"D4",x"AA",x"68",x"13",x"6D",x"96",x"DA",x"2A", -- 0x0708
		x"B5",x"AB",x"43",x"5B",x"87",x"A7",x"57",x"57", -- 0x0710
		x"8F",x"8F",x"1F",x"3F",x"7F",x"7F",x"FB",x"FF", -- 0x0718
		x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"E7",x"A3", -- 0x0720
		x"F2",x"51",x"75",x"4B",x"2E",x"38",x"45",x"71", -- 0x0728
		x"F8",x"FC",x"FE",x"FF",x"FC",x"FE",x"F8",x"89", -- 0x0730
		x"C8",x"84",x"06",x"A4",x"9D",x"42",x"B4",x"58", -- 0x0738
		x"D4",x"98",x"EA",x"D5",x"59",x"76",x"23",x"B7", -- 0x0740
		x"9F",x"C7",x"DF",x"FF",x"FF",x"FB",x"FF",x"FF", -- 0x0748
		x"08",x"54",x"84",x"48",x"AD",x"7A",x"50",x"21", -- 0x0750
		x"F4",x"68",x"3C",x"8F",x"E3",x"FA",x"FC",x"F8", -- 0x0758
		x"D1",x"20",x"A8",x"F5",x"2F",x"9F",x"8F",x"DF", -- 0x0760
		x"2F",x"C7",x"E7",x"FF",x"7F",x"1F",x"3F",x"1F", -- 0x0768
		x"47",x"D1",x"6D",x"1F",x"CF",x"FE",x"FF",x"BF", -- 0x0770
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"FD",x"FF", -- 0x0778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0788
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0790
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F8
		x"FF",x"33",x"21",x"59",x"8E",x"62",x"7F",x"FF", -- 0x0800
		x"7F",x"7F",x"7F",x"03",x"03",x"F3",x"F3",x"F3", -- 0x0808
		x"FF",x"C7",x"03",x"AB",x"D3",x"77",x"0F",x"D7", -- 0x0810
		x"C7",x"F3",x"C3",x"E9",x"E9",x"F7",x"C3",x"F3", -- 0x0818
		x"F3",x"F3",x"F3",x"F3",x"F3",x"F0",x"F1",x"FF", -- 0x0820
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"B0", -- 0x0828
		x"E3",x"C9",x"F3",x"C3",x"87",x"D3",x"67",x"47", -- 0x0830
		x"2F",x"83",x"E3",x"81",x"81",x"53",x"27",x"A3", -- 0x0838
		x"00",x"54",x"47",x"D3",x"8F",x"C6",x"73",x"0F", -- 0x0840
		x"E7",x"E7",x"15",x"A3",x"93",x"C4",x"F8",x"0D", -- 0x0848
		x"17",x"03",x"8F",x"C7",x"9F",x"5F",x"7F",x"FF", -- 0x0850
		x"E7",x"A3",x"D3",x"71",x"61",x"2B",x"93",x"C7", -- 0x0858
		x"10",x"88",x"98",x"0D",x"0F",x"05",x"40",x"20", -- 0x0860
		x"06",x"0C",x"C6",x"E3",x"D0",x"4E",x"FF",x"FF", -- 0x0868
		x"2F",x"BF",x"1F",x"9F",x"8F",x"0F",x"47",x"DF", -- 0x0870
		x"67",x"67",x"DF",x"9F",x"DF",x"3F",x"FF",x"FF", -- 0x0878
		x"FF",x"F1",x"C8",x"C9",x"47",x"A8",x"10",x"09", -- 0x0880
		x"11",x"58",x"AC",x"9D",x"EE",x"F2",x"F9",x"99", -- 0x0888
		x"FF",x"9F",x"D7",x"C3",x"A3",x"C3",x"2B",x"15", -- 0x0890
		x"01",x"89",x"89",x"05",x"97",x"23",x"1F",x"1F", -- 0x0898
		x"E0",x"92",x"DA",x"CB",x"ED",x"FD",x"C8",x"E8", -- 0x08A0
		x"F0",x"F8",x"E8",x"6E",x"B4",x"8D",x"86",x"40", -- 0x08A8
		x"1F",x"87",x"C3",x"D3",x"6F",x"FF",x"6F",x"3F", -- 0x08B0
		x"3F",x"A7",x"C3",x"23",x"A9",x"19",x"13",x"0D", -- 0x08B8
		x"20",x"C1",x"C8",x"39",x"9F",x"18",x"10",x"89", -- 0x08C0
		x"91",x"D8",x"AC",x"5D",x"4E",x"E2",x"E9",x"F1", -- 0x08C8
		x"A3",x"9B",x"D7",x"DF",x"AF",x"CF",x"23",x"11", -- 0x08D0
		x"01",x"89",x"9F",x"2F",x"9F",x"27",x"21",x"19", -- 0x08D8
		x"A0",x"9A",x"CE",x"B3",x"8D",x"D5",x"88",x"40", -- 0x08E0
		x"71",x"38",x"88",x"EE",x"F7",x"F7",x"FF",x"FF", -- 0x08E8
		x"11",x"A1",x"E3",x"D7",x"3F",x"0F",x"3F",x"0F", -- 0x08F0
		x"03",x"21",x"C1",x"6F",x"3F",x"9F",x"FF",x"FF", -- 0x08F8
		x"FF",x"F9",x"F9",x"D0",x"CB",x"F7",x"C7",x"EF", -- 0x0900
		x"E7",x"D2",x"E0",x"B0",x"80",x"CB",x"E3",x"D7", -- 0x0908
		x"FF",x"F3",x"E1",x"E8",x"9A",x"ED",x"FF",x"FF", -- 0x0910
		x"7F",x"7E",x"7E",x"06",x"0E",x"FF",x"FF",x"FF", -- 0x0918
		x"83",x"C0",x"ED",x"C7",x"97",x"C7",x"A3",x"A1", -- 0x0920
		x"81",x"95",x"C9",x"E3",x"D3",x"C0",x"F0",x"D4", -- 0x0928
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0930
		x"FF",x"FB",x"F3",x"C9",x"A1",x"9D",x"C2",x"68", -- 0x0938
		x"C8",x"E7",x"F3",x"FE",x"FF",x"E9",x"B0",x"A2", -- 0x0940
		x"B7",x"80",x"D4",x"F0",x"B8",x"94",x"DD",x"FE", -- 0x0948
		x"E4",x"A0",x"16",x"9A",x"2F",x"8D",x"DC",x"52", -- 0x0950
		x"B1",x"F1",x"41",x"A8",x"30",x"1C",x"25",x"77", -- 0x0958
		x"F8",x"EA",x"ED",x"EA",x"F4",x"D6",x"DA",x"DB", -- 0x0960
		x"ED",x"F6",x"F5",x"EE",x"E7",x"F1",x"FF",x"FF", -- 0x0968
		x"27",x"42",x"E1",x"88",x"10",x"5D",x"82",x"62", -- 0x0970
		x"B0",x"5A",x"64",x"BD",x"9F",x"DD",x"C7",x"FF", -- 0x0978
		x"FF",x"FC",x"F8",x"E9",x"E7",x"F0",x"F0",x"E9", -- 0x0980
		x"D1",x"D0",x"D8",x"CD",x"E2",x"FA",x"FE",x"F3", -- 0x0988
		x"FF",x"FB",x"75",x"01",x"90",x"CA",x"28",x"14", -- 0x0990
		x"00",x"88",x"8A",x"07",x"21",x"97",x"4F",x"FF", -- 0x0998
		x"F8",x"F0",x"D4",x"C8",x"ED",x"E7",x"F0",x"FC", -- 0x09A0
		x"F6",x"F5",x"F9",x"EF",x"E1",x"F1",x"E8",x"F0", -- 0x09A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x09B0
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FF", -- 0x09B8
		x"C8",x"ED",x"E7",x"F7",x"FF",x"FD",x"F8",x"E8", -- 0x09C0
		x"EB",x"E5",x"F1",x"F8",x"F4",x"F6",x"F8",x"E8", -- 0x09C8
		x"FD",x"FD",x"FC",x"FE",x"FF",x"FF",x"FF",x"FD", -- 0x09D0
		x"FD",x"FC",x"FE",x"FE",x"7F",x"7F",x"FF",x"FF", -- 0x09D8
		x"E1",x"F5",x"F0",x"EA",x"EC",x"E3",x"FB",x"FF", -- 0x09E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FA",x"F8", -- 0x09F0
		x"F0",x"DA",x"C5",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x09F8
		x"FF",x"FF",x"FF",x"DF",x"DF",x"C0",x"FF",x"EF", -- 0x0A00
		x"CF",x"CF",x"C3",x"C7",x"FF",x"DF",x"DF",x"DF", -- 0x0A08
		x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F0",x"F0", -- 0x0A10
		x"E0",x"E0",x"C0",x"C0",x"81",x"81",x"83",x"83", -- 0x0A18
		x"C7",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC", -- 0x0A20
		x"FC",x"FC",x"FC",x"F8",x"F8",x"FF",x"FF",x"F8", -- 0x0A28
		x"07",x"07",x"0F",x"0F",x"07",x"07",x"07",x"17", -- 0x0A30
		x"11",x"1F",x"0F",x"0F",x"07",x"FF",x"FF",x"3F", -- 0x0A38
		x"F0",x"F0",x"F0",x"F0",x"F0",x"E0",x"E0",x"E0", -- 0x0A40
		x"E0",x"C0",x"C0",x"C1",x"C1",x"81",x"83",x"83", -- 0x0A48
		x"3F",x"6F",x"6F",x"6F",x"63",x"7F",x"EF",x"EF", -- 0x0A50
		x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"E3",x"FF", -- 0x0A58
		x"03",x"07",x"07",x"07",x"0F",x"1F",x"3F",x"3B", -- 0x0A60
		x"7B",x"7B",x"D8",x"DF",x"DF",x"C0",x"FF",x"FF", -- 0x0A68
		x"DF",x"C7",x"FF",x"FF",x"FF",x"DF",x"9F",x"9F", -- 0x0A70
		x"9F",x"9F",x"9F",x"DF",x"C3",x"07",x"FF",x"FF", -- 0x0A78
		x"00",x"3F",x"3F",x"3E",x"20",x"01",x"0F",x"3F", -- 0x0A80
		x"3F",x"3F",x"30",x"21",x"3F",x"3F",x"3F",x"26", -- 0x0A88
		x"00",x"F8",x"C0",x"06",x"3E",x"FE",x"FE",x"FE", -- 0x0A90
		x"FE",x"E2",x"FE",x"FE",x"FE",x"FE",x"F2",x"7E", -- 0x0A98
		x"3F",x"1F",x"03",x"3F",x"3F",x"3F",x"3F",x"33", -- 0x0AA0
		x"27",x"00",x"00",x"3F",x"3F",x"3E",x"3E",x"33", -- 0x0AA8
		x"FE",x"FE",x"FE",x"FE",x"1A",x"FE",x"DE",x"DE", -- 0x0AB0
		x"42",x"00",x"00",x"FE",x"FE",x"1E",x"3E",x"FE", -- 0x0AB8
		x"27",x"3E",x"3C",x"3C",x"3C",x"3C",x"27",x"03", -- 0x0AC0
		x"01",x"38",x"3F",x"3F",x"3F",x"3E",x"3E",x"3E", -- 0x0AC8
		x"F2",x"06",x"0E",x"0E",x"0E",x"1E",x"FE",x"FE", -- 0x0AD0
		x"3E",x"0A",x"1E",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0AD8
		x"3E",x"22",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x0AE0
		x"30",x"21",x"3F",x"3F",x"3F",x"38",x"00",x"00", -- 0x0AE8
		x"E2",x"7E",x"FE",x"FE",x"C6",x"FE",x"DE",x"C2", -- 0x0AF0
		x"FE",x"FE",x"FE",x"FE",x"FE",x"E2",x"00",x"00", -- 0x0AF8
		x"00",x"3F",x"77",x"71",x"7F",x"77",x"77",x"51", -- 0x0B00
		x"00",x"00",x"00",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x0B08
		x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"C2",x"86", -- 0x0B10
		x"00",x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0B18
		x"27",x"3E",x"3F",x"3E",x"3E",x"3E",x"32",x"26", -- 0x0B20
		x"3F",x"3F",x"3F",x"3F",x"3F",x"31",x"23",x"3F", -- 0x0B28
		x"02",x"1E",x"FE",x"FE",x"E2",x"FE",x"DE",x"42", -- 0x0B30
		x"FE",x"FE",x"FE",x"FE",x"FE",x"C2",x"86",x"FE", -- 0x0B38
		x"3F",x"3F",x"3C",x"3D",x"3F",x"3D",x"3D",x"3C", -- 0x0B40
		x"27",x"08",x"00",x"03",x"3F",x"3F",x"3F",x"31", -- 0x0B48
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"C2",x"80", -- 0x0B50
		x"00",x"0E",x"7E",x"FE",x"7E",x"7E",x"7E",x"3E", -- 0x0B58
		x"23",x"3F",x"3F",x"3F",x"3F",x"21",x"3F",x"3F", -- 0x0B60
		x"3F",x"3F",x"3F",x"3F",x"30",x"21",x"00",x"00", -- 0x0B68
		x"F2",x"FE",x"EE",x"EE",x"E2",x"BE",x"FE",x"FE", -- 0x0B70
		x"FE",x"FE",x"FE",x"FE",x"E2",x"C6",x"00",x"00", -- 0x0B78
		x"FF",x"FF",x"FF",x"DF",x"DE",x"DE",x"DF",x"DF", -- 0x0B80
		x"C3",x"FF",x"DF",x"DF",x"DF",x"C1",x"FF",x"FF", -- 0x0B88
		x"FF",x"E7",x"87",x"83",x"C3",x"21",x"A9",x"9B", -- 0x0B90
		x"E7",x"A3",x"93",x"D9",x"C1",x"63",x"27",x"FF", -- 0x0B98
		x"00",x"3F",x"3B",x"3B",x"3B",x"3B",x"3B",x"20", -- 0x0BA0
		x"3F",x"3F",x"3E",x"3E",x"23",x"3F",x"3F",x"3F", -- 0x0BA8
		x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"C2", -- 0x0BB0
		x"86",x"E0",x"C0",x"40",x"C0",x"C0",x"C0",x"C0", -- 0x0BB8
		x"3F",x"27",x"3F",x"3F",x"3F",x"3F",x"3F",x"31", -- 0x0BC0
		x"23",x"30",x"00",x"0F",x"3F",x"3F",x"3F",x"33", -- 0x0BC8
		x"C2",x"7E",x"F6",x"F6",x"F6",x"F6",x"F2",x"9E", -- 0x0BD0
		x"E0",x"00",x"0E",x"FE",x"FE",x"FE",x"F2",x"FE", -- 0x0BD8
		x"27",x"3F",x"1F",x"1F",x"1E",x"02",x"3F",x"3F", -- 0x0BE0
		x"3F",x"3F",x"3F",x"3F",x"30",x"21",x"00",x"00", -- 0x0BE8
		x"FE",x"3E",x"FE",x"FE",x"FE",x"32",x"FE",x"FE", -- 0x0BF0
		x"FE",x"FE",x"FE",x"FE",x"E2",x"C6",x"00",x"00", -- 0x0BF8
		x"00",x"F3",x"E7",x"E7",x"CF",x"CC",x"9F",x"BE", -- 0x0C00
		x"3E",x"3E",x"7F",x"62",x"7E",x"7E",x"43",x"7F", -- 0x0C08
		x"00",x"FE",x"FE",x"FE",x"FE",x"72",x"E6",x"FE", -- 0x0C10
		x"FE",x"7E",x"E2",x"FE",x"FE",x"62",x"FE",x"FE", -- 0x0C18
		x"7F",x"6D",x"00",x"00",x"7F",x"7F",x"7F",x"7F", -- 0x0C20
		x"5F",x"7F",x"7C",x"79",x"7F",x"5F",x"00",x"00", -- 0x0C28
		x"FE",x"FE",x"80",x"00",x"FE",x"FE",x"FE",x"FE", -- 0x0C30
		x"CE",x"9E",x"FE",x"FE",x"FA",x"F6",x"80",x"00", -- 0x0C38
		x"00",x"FE",x"FC",x"FC",x"FC",x"07",x"FF",x"DF", -- 0x0C40
		x"DF",x"DF",x"C2",x"70",x"81",x"0F",x"7F",x"FF", -- 0x0C48
		x"00",x"0E",x"0E",x"06",x"16",x"FA",x"FE",x"FE", -- 0x0C50
		x"88",x"00",x"06",x"3E",x"FE",x"EE",x"EE",x"E6", -- 0x0C58
		x"FF",x"FF",x"F1",x"FF",x"1D",x"E4",x"FF",x"FF", -- 0x0C60
		x"FF",x"BF",x"FF",x"FF",x"FC",x"38",x"00",x"00", -- 0x0C68
		x"3E",x"FE",x"FE",x"FE",x"FE",x"62",x"FE",x"FE", -- 0x0C70
		x"FA",x"FE",x"EE",x"EE",x"6E",x"E2",x"00",x"00", -- 0x0C78
		x"00",x"FE",x"FE",x"FC",x"FC",x"FC",x"39",x"78", -- 0x0C80
		x"00",x"03",x"F3",x"F3",x"E7",x"E6",x"00",x"00", -- 0x0C88
		x"00",x"7E",x"F6",x"F6",x"F6",x"82",x"FE",x"EE", -- 0x0C90
		x"22",x"FE",x"FE",x"FE",x"FE",x"C2",x"00",x"00", -- 0x0C98
		x"00",x"FF",x"F7",x"F1",x"FF",x"1F",x"FF",x"FF", -- 0x0CA0
		x"FF",x"F8",x"F1",x"FF",x"37",x"70",x"00",x"00", -- 0x0CA8
		x"00",x"FE",x"FE",x"FE",x"FE",x"C2",x"E0",x"C0", -- 0x0CB0
		x"C0",x"C0",x"C0",x"C6",x"FE",x"FE",x"00",x"00", -- 0x0CB8
		x"FF",x"FF",x"FF",x"EF",x"EF",x"EF",x"E3",x"FF", -- 0x0CC0
		x"1E",x"E4",x"60",x"4C",x"68",x"3C",x"83",x"F0", -- 0x0CC8
		x"FF",x"E7",x"C3",x"A1",x"41",x"53",x"5B",x"E1", -- 0x0CD0
		x"B1",x"E1",x"75",x"1F",x"07",x"BF",x"FF",x"FF", -- 0x0CD8
		x"00",x"FF",x"FF",x"FF",x"FF",x"F0",x"FF",x"3F", -- 0x0CE0
		x"3F",x"3F",x"32",x"3E",x"3E",x"62",x"00",x"00", -- 0x0CE8
		x"00",x"FE",x"FE",x"FE",x"FE",x"C2",x"FE",x"EE", -- 0x0CF0
		x"22",x"FE",x"FE",x"FE",x"FE",x"62",x"00",x"00", -- 0x0CF8
		x"00",x"3F",x"3F",x"3F",x"3F",x"3F",x"30",x"20", -- 0x0D00
		x"00",x"00",x"3F",x"3F",x"3E",x"3E",x"3E",x"22", -- 0x0D08
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"01", -- 0x0D10
		x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F", -- 0x0D18
		x"3F",x"3F",x"3F",x"3F",x"3E",x"27",x"3F",x"3F", -- 0x0D20
		x"3F",x"27",x"3F",x"3F",x"3F",x"26",x"00",x"00", -- 0x0D28
		x"F9",x"FF",x"F0",x"E0",x"20",x"E0",x"E0",x"E0", -- 0x0D30
		x"E1",x"FF",x"FF",x"F1",x"3F",x"7F",x"10",x"00", -- 0x0D38
		x"00",x"3F",x"3F",x"3F",x"3F",x"21",x"3F",x"3F", -- 0x0D40
		x"3E",x"3E",x"23",x"3F",x"1F",x"1F",x"1F",x"03", -- 0x0D48
		x"00",x"FF",x"FF",x"FF",x"FF",x"C7",x"8F",x"FF", -- 0x0D50
		x"FF",x"1F",x"FF",x"F8",x"FF",x"FC",x"00",x"03", -- 0x0D58
		x"38",x"03",x"07",x"3F",x"3F",x"26",x"04",x"07", -- 0x0D60
		x"05",x"04",x"07",x"00",x"00",x"02",x"00",x"00", -- 0x0D68
		x"07",x"F7",x"F7",x"F7",x"F4",x"17",x"33",x"F3", -- 0x0D70
		x"F3",x"31",x"F7",x"F7",x"F7",x"F4",x"00",x"00", -- 0x0D78
		x"00",x"3F",x"3F",x"3F",x"3F",x"30",x"3F",x"3B", -- 0x0D80
		x"3B",x"3B",x"38",x"3F",x"3D",x"24",x"00",x"00", -- 0x0D88
		x"00",x"9F",x"9F",x"9F",x"9F",x"9F",x"98",x"90", -- 0x0D90
		x"80",x"80",x"9F",x"97",x"97",x"90",x"00",x"00", -- 0x0D98
		x"00",x"3F",x"1F",x"07",x"3F",x"3F",x"3F",x"3F", -- 0x0DA0
		x"26",x"3F",x"2F",x"23",x"3F",x"3F",x"20",x"00", -- 0x0DA8
		x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"EB",x"EF", -- 0x0DB0
		x"2F",x"EF",x"EF",x"EF",x"EC",x"28",x"00",x"00", -- 0x0DB8
		x"00",x"3F",x"1F",x"01",x"3F",x"3F",x"27",x"3F", -- 0x0DC0
		x"1F",x"1F",x"0F",x"3F",x"3E",x"2C",x"00",x"00", -- 0x0DC8
		x"00",x"FF",x"FF",x"FE",x"FE",x"86",x"FE",x"FE", -- 0x0DD0
		x"FE",x"FF",x"FF",x"FF",x"63",x"FF",x"00",x"00", -- 0x0DD8
		x"00",x"3F",x"3F",x"3F",x"3B",x"3B",x"2B",x"3B", -- 0x0DE0
		x"18",x"0F",x"3F",x"3F",x"38",x"30",x"00",x"00", -- 0x0DE8
		x"00",x"3F",x"8F",x"8D",x"C5",x"CD",x"E5",x"E4", -- 0x0DF0
		x"F3",x"F3",x"F9",x"F9",x"1D",x"3D",x"00",x"00", -- 0x0DF8
		x"00",x"3F",x"3F",x"3F",x"3C",x"38",x"3F",x"2F", -- 0x0E00
		x"04",x"00",x"3F",x"2D",x"2D",x"8D",x"C4",x"E7", -- 0x0E08
		x"00",x"FE",x"F6",x"F6",x"16",x"32",x"FE",x"FE", -- 0x0E10
		x"80",x"00",x"FE",x"FE",x"F6",x"F6",x"16",x"06", -- 0x0E18
		x"FE",x"FE",x"E2",x"A3",x"A7",x"B1",x"99",x"D1", -- 0x0E20
		x"C7",x"F1",x"FA",x"FA",x"FB",x"F8",x"FE",x"FF", -- 0x0E28
		x"F3",x"FF",x"17",x"F7",x"F7",x"F3",x"FF",x"7F", -- 0x0E30
		x"3F",x"2F",x"07",x"87",x"53",x"A7",x"2F",x"FF", -- 0x0E38
		x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"C4", -- 0x0E40
		x"8C",x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"FC", -- 0x0E48
		x"00",x"FE",x"FE",x"FE",x"FE",x"86",x"FE",x"FE", -- 0x0E50
		x"FE",x"FE",x"7E",x"E2",x"90",x"00",x"7E",x"FE", -- 0x0E58
		x"FC",x"E4",x"CC",x"FC",x"FC",x"FC",x"FC",x"F5", -- 0x0E60
		x"3D",x"FD",x"FD",x"FD",x"FD",x"84",x"00",x"00", -- 0x0E68
		x"FE",x"86",x"FE",x"FE",x"FE",x"7E",x"E2",x"FE", -- 0x0E70
		x"FE",x"FE",x"FE",x"FE",x"7E",x"E6",x"00",x"00", -- 0x0E78
		x"00",x"3F",x"3F",x"3F",x"3F",x"3F",x"2F",x"3E", -- 0x0E80
		x"3F",x"3F",x"3F",x"3F",x"3F",x"31",x"23",x"3F", -- 0x0E88
		x"00",x"FE",x"FE",x"86",x"8E",x"FE",x"FE",x"F2", -- 0x0E90
		x"E6",x"FE",x"FE",x"FE",x"C6",x"FE",x"FE",x"FE", -- 0x0E98
		x"1F",x"1F",x"1F",x"07",x"3F",x"3F",x"1E",x"3F", -- 0x0EA0
		x"3F",x"3F",x"3F",x"3F",x"20",x"3F",x"00",x"00", -- 0x0EA8
		x"FE",x"FE",x"F2",x"FE",x"EE",x"2E",x"66",x"FE", -- 0x0EB0
		x"FE",x"FE",x"FE",x"FE",x"62",x"FE",x"00",x"00", -- 0x0EB8
		x"00",x"3F",x"3F",x"3F",x"21",x"3F",x"3F",x"3D", -- 0x0EC0
		x"3D",x"24",x"3F",x"3F",x"3F",x"3F",x"38",x"00", -- 0x0EC8
		x"00",x"FE",x"FE",x"FE",x"86",x"06",x"F6",x"F6", -- 0x0ED0
		x"F2",x"1E",x"FE",x"FE",x"FE",x"FE",x"66",x"40", -- 0x0ED8
		x"00",x"3F",x"7F",x"7F",x"7F",x"7F",x"7E",x"5C", -- 0x0EE0
		x"3F",x"3F",x"23",x"3F",x"1F",x"03",x"00",x"00", -- 0x0EE8
		x"00",x"FE",x"F6",x"F6",x"F6",x"F6",x"12",x"3E", -- 0x0EF0
		x"FE",x"FE",x"FE",x"FE",x"FE",x"62",x"00",x"00", -- 0x0EF8
		x"00",x"3F",x"3E",x"22",x"3E",x"3F",x"3F",x"3F", -- 0x0F00
		x"3F",x"23",x"00",x"00",x"3F",x"3F",x"2F",x"2F", -- 0x0F08
		x"00",x"FF",x"FF",x"FF",x"31",x"FF",x"FF",x"FF", -- 0x0F10
		x"C1",x"83",x"00",x"00",x"FF",x"FF",x"FF",x"E7", -- 0x0F18
		x"20",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3E", -- 0x0F20
		x"3E",x"3F",x"3F",x"3F",x"30",x"20",x"00",x"00", -- 0x0F28
		x"FF",x"FF",x"FF",x"FF",x"F9",x"1F",x"F7",x"F7", -- 0x0F30
		x"17",x"F7",x"F1",x"FF",x"1F",x"39",x"00",x"00", -- 0x0F38
		x"FF",x"F5",x"F0",x"D8",x"A0",x"B4",x"99",x"C7", -- 0x0F40
		x"F3",x"FF",x"FF",x"FF",x"DF",x"DE",x"DE",x"C2", -- 0x0F48
		x"FF",x"FF",x"EF",x"6F",x"6F",x"E1",x"FF",x"DF", -- 0x0F50
		x"C7",x"FF",x"FF",x"FF",x"FF",x"F7",x"F7",x"F0", -- 0x0F58
		x"3E",x"3E",x"3E",x"3F",x"23",x"3F",x"3F",x"3F", -- 0x0F60
		x"3F",x"30",x"21",x"3F",x"2F",x"23",x"00",x"00", -- 0x0F68
		x"FF",x"FB",x"1B",x"F8",x"FF",x"FF",x"FF",x"CF", -- 0x0F70
		x"9C",x"87",x"07",x"07",x"07",x"0D",x"00",x"00", -- 0x0F78
		x"00",x"3F",x"3F",x"3F",x"3F",x"30",x"20",x"3F", -- 0x0F80
		x"3F",x"3F",x"27",x"3F",x"3F",x"3F",x"3C",x"2F", -- 0x0F88
		x"00",x"FE",x"DE",x"DE",x"DE",x"42",x"FE",x"FE", -- 0x0F90
		x"FE",x"86",x"FE",x"FE",x"FE",x"FE",x"1E",x"FA", -- 0x0F98
		x"3B",x"1B",x"08",x"3F",x"3F",x"3F",x"3F",x"30", -- 0x0FA0
		x"3F",x"3F",x"3F",x"3F",x"30",x"20",x"00",x"00", -- 0x0FA8
		x"C0",x"80",x"80",x"80",x"82",x"FE",x"FE",x"FE", -- 0x0FB0
		x"FE",x"FE",x"E2",x"FE",x"5E",x"C2",x"00",x"00", -- 0x0FB8
		x"00",x"3F",x"3F",x"3F",x"3F",x"3C",x"21",x"0E", -- 0x0FC0
		x"00",x"00",x"3F",x"1F",x"1F",x"07",x"3F",x"3F", -- 0x0FC8
		x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"32",x"66", -- 0x0FD0
		x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"82",x"06", -- 0x0FD8
		x"3F",x"27",x"0F",x"07",x"22",x"31",x"38",x"1C", -- 0x0FE0
		x"1E",x"1F",x"1F",x"0F",x"3F",x"3C",x"00",x"00", -- 0x0FE8
		x"FE",x"FE",x"FE",x"F2",x"3E",x"FE",x"FE",x"7E", -- 0x0FF0
		x"22",x"9E",x"86",x"C2",x"E2",x"F0",x"00",x"00", -- 0x0FF8
		x"00",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"23", -- 0x1000
		x"3F",x"00",x"00",x"3F",x"3D",x"3D",x"3C",x"00", -- 0x1008
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"46",x"60", -- 0x1010
		x"6F",x"6F",x"6F",x"E7",x"E7",x"E7",x"03",x"1F", -- 0x1018
		x"00",x"3C",x"3C",x"3C",x"3C",x"24",x"00",x"00", -- 0x1020
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"31",x"3F", -- 0x1028
		x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"EE",x"60", -- 0x1030
		x"0E",x"9E",x"DE",x"D6",x"D6",x"D6",x"D2",x"C0", -- 0x1038
		x"01",x"3C",x"3F",x"3F",x"3F",x"23",x"00",x"00", -- 0x1040
		x"3E",x"3E",x"3E",x"3E",x"3E",x"26",x"3E",x"00", -- 0x1048
		x"FF",x"7F",x"7F",x"73",x"7B",x"7B",x"7B",x"00", -- 0x1050
		x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"40",x"7F", -- 0x1058
		x"00",x"3F",x"3F",x"3F",x"3F",x"3F",x"21",x"3F", -- 0x1060
		x"38",x"38",x"39",x"39",x"39",x"29",x"00",x"00", -- 0x1068
		x"00",x"3E",x"3E",x"3E",x"3E",x"3E",x"36",x"3E", -- 0x1070
		x"3E",x"3C",x"FD",x"F9",x"F3",x"E7",x"07",x"03", -- 0x1078
		x"C0",x"DC",x"DC",x"DC",x"CC",x"E6",x"EE",x"EE", -- 0x1080
		x"EE",x"6E",x"62",x"7E",x"3E",x"7E",x"72",x"00", -- 0x1088
		x"00",x"FC",x"F8",x"F9",x"FB",x"83",x"E7",x"E7", -- 0x1090
		x"07",x"07",x"FF",x"FF",x"FF",x"C7",x"F7",x"07", -- 0x1098
		x"00",x"3C",x"1C",x"1C",x"1C",x"0C",x"00",x"80", -- 0x10A0
		x"9F",x"9F",x"BF",x"BF",x"BF",x"B0",x"BE",x"80", -- 0x10A8
		x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"82",x"00", -- 0x10B0
		x"BF",x"BF",x"00",x"00",x"FE",x"7E",x"7E",x"00", -- 0x10B8
		x"00",x"7B",x"7B",x"79",x"7D",x"7C",x"5D",x"01", -- 0x10C0
		x"BD",x"BD",x"BD",x"BD",x"BD",x"B5",x"80",x"00", -- 0x10C8
		x"03",x"FB",x"FB",x"FB",x"3B",x"03",x"FF",x"FF", -- 0x10D0
		x"E0",x"FE",x"FE",x"FE",x"FE",x"06",x"00",x"00", -- 0x10D8
		x"80",x"BF",x"BF",x"9F",x"9F",x"9F",x"87",x"00", -- 0x10E0
		x"00",x"7E",x"7E",x"7E",x"7E",x"46",x"00",x"00", -- 0x10E8
		x"03",x"7B",x"7B",x"7B",x"49",x"7D",x"7D",x"01", -- 0x10F0
		x"FC",x"FE",x"FE",x"FE",x"FE",x"CE",x"00",x"00", -- 0x10F8
		x"C0",x"DF",x"DF",x"D1",x"C0",x"00",x"7F",x"FE", -- 0x1100
		x"FC",x"FC",x"FD",x"8D",x"7D",x"7D",x"00",x"00", -- 0x1108
		x"00",x"F8",x"F2",x"E6",x"0E",x"1E",x"3E",x"72", -- 0x1110
		x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"80",x"00", -- 0x1118
		x"FC",x"01",x"01",x"7F",x"7F",x"7F",x"7C",x"78", -- 0x1120
		x"78",x"01",x"01",x"79",x"79",x"79",x"78",x"00", -- 0x1128
		x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"4E",x"0A", -- 0x1130
		x"0E",x"FE",x"FE",x"FE",x"FE",x"C6",x"00",x"00", -- 0x1138
		x"E0",x"FF",x"FF",x"78",x"78",x"7C",x"4D",x"7D", -- 0x1140
		x"7D",x"7D",x"7D",x"7D",x"3D",x"0D",x"01",x"01", -- 0x1148
		x"00",x"FC",x"FC",x"FC",x"8C",x"1C",x"80",x"80", -- 0x1150
		x"9C",x"9C",x"9C",x"9C",x"9C",x"94",x"80",x"80", -- 0x1158
		x"03",x"7B",x"7A",x"78",x"78",x"79",x"79",x"59", -- 0x1160
		x"00",x"00",x"7D",x"7D",x"7D",x"7D",x"65",x"01", -- 0x1168
		x"80",x"3C",x"3C",x"7C",x"FC",x"FC",x"FC",x"CC", -- 0x1170
		x"00",x"00",x"FC",x"FC",x"E4",x"E4",x"E0",x"F0", -- 0x1178
		x"FF",x"00",x"00",x"DF",x"DF",x"DF",x"DF",x"DF", -- 0x1180
		x"D3",x"DF",x"DF",x"C1",x"C1",x"FD",x"FD",x"FD", -- 0x1188
		x"FF",x"1F",x"1F",x"DB",x"DF",x"DF",x"DF",x"DF", -- 0x1190
		x"DF",x"FF",x"F8",x"F8",x"0F",x"FF",x"FF",x"FF", -- 0x1198
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x11A0
		x"FF",x"FB",x"FB",x"F8",x"FF",x"FF",x"FF",x"FF", -- 0x11A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11B0
		x"EF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x11B8
		x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF", -- 0x11C0
		x"E9",x"00",x"00",x"FD",x"ED",x"FD",x"FD",x"FD", -- 0x11C8
		x"FF",x"FF",x"FF",x"FF",x"20",x"7F",x"7F",x"7F", -- 0x11D0
		x"7F",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11D8
		x"FD",x"FD",x"FD",x"FD",x"FD",x"C5",x"00",x"00", -- 0x11E0
		x"DF",x"DF",x"DF",x"DF",x"DF",x"DF",x"CF",x"C0", -- 0x11E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"0B", -- 0x11F0
		x"E0",x"E0",x"FF",x"FF",x"3F",x"77",x"7F",x"7F", -- 0x11F8
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"03", -- 0x1200
		x"FD",x"DE",x"FF",x"FE",x"FA",x"F5",x"E8",x"E8", -- 0x1208
		x"FF",x"9F",x"5B",x"A5",x"E5",x"C1",x"6B",x"3F", -- 0x1210
		x"8F",x"EF",x"FF",x"FF",x"3F",x"FF",x"FF",x"BF", -- 0x1218
		x"ED",x"F3",x"D2",x"CD",x"E9",x"E4",x"F6",x"F0", -- 0x1220
		x"F0",x"EC",x"E9",x"ED",x"E5",x"33",x"C3",x"8F", -- 0x1228
		x"BF",x"BF",x"3F",x"0F",x"FF",x"FF",x"FF",x"3F", -- 0x1230
		x"BF",x"BF",x"BF",x"BF",x"BF",x"87",x"FF",x"FF", -- 0x1238
		x"A7",x"C3",x"0B",x"58",x"FF",x"BF",x"3F",x"FF", -- 0x1240
		x"DF",x"DF",x"DF",x"DF",x"FF",x"FF",x"FF",x"07", -- 0x1248
		x"FF",x"FF",x"FF",x"1F",x"DF",x"DF",x"DF",x"DF", -- 0x1250
		x"DF",x"DF",x"DF",x"DF",x"DF",x"DF",x"C7",x"FF", -- 0x1258
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"7E", -- 0x1260
		x"38",x"8A",x"1C",x"DF",x"4D",x"E7",x"FF",x"FF", -- 0x1268
		x"FF",x"E7",x"C7",x"A3",x"E3",x"4B",x"71",x"21", -- 0x1270
		x"B1",x"63",x"EB",x"6B",x"37",x"9F",x"FF",x"FF", -- 0x1278
		x"61",x"3F",x"9F",x"FF",x"7F",x"FF",x"FF",x"E0", -- 0x1280
		x"FF",x"FC",x"FE",x"FC",x"EC",x"2E",x"E7",x"F3", -- 0x1288
		x"80",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"00", -- 0x1290
		x"FF",x"7C",x"08",x"38",x"16",x"88",x"11",x"A1", -- 0x1298
		x"FB",x"F8",x"FC",x"E5",x"FD",x"FC",x"F8",x"EE", -- 0x12A0
		x"35",x"F3",x"A3",x"B9",x"8C",x"E6",x"FF",x"FF", -- 0x12A8
		x"60",x"32",x"AF",x"97",x"4E",x"80",x"00",x"20", -- 0x12B0
		x"A4",x"14",x"2C",x"DF",x"D1",x"24",x"98",x"CC", -- 0x12B8
		x"FF",x"E0",x"FF",x"FF",x"F8",x"F5",x"F4",x"FF", -- 0x12C0
		x"EF",x"EA",x"E2",x"37",x"F3",x"CA",x"A4",x"83", -- 0x12C8
		x"FA",x"62",x"A6",x"F3",x"41",x"61",x"A1",x"F3", -- 0x12D0
		x"43",x"67",x"07",x"15",x"18",x"A9",x"64",x"6E", -- 0x12D8
		x"48",x"D0",x"F8",x"F5",x"6B",x"0F",x"FF",x"FF", -- 0x12E0
		x"1E",x"21",x"09",x"D0",x"7C",x"39",x"8F",x"E7", -- 0x12E8
		x"74",x"37",x"99",x"CF",x"FF",x"FF",x"F8",x"C1", -- 0x12F0
		x"30",x"F8",x"F8",x"D0",x"6A",x"37",x"9F",x"FF", -- 0x12F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"00", -- 0x1300
		x"FF",x"FF",x"63",x"21",x"11",x"81",x"05",x"AB", -- 0x1308
		x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"7F",x"00", -- 0x1310
		x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"00",x"FE", -- 0x1318
		x"C7",x"6F",x"20",x"C0",x"40",x"41",x"7F",x"7F", -- 0x1320
		x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"CF",x"8F", -- 0x1328
		x"FE",x"FE",x"CE",x"8E",x"8E",x"8E",x"86",x"06", -- 0x1330
		x"06",x"06",x"06",x"06",x"06",x"0E",x"8F",x"8F", -- 0x1338
		x"80",x"00",x"00",x"7C",x"FA",x"F4",x"DD",x"C6", -- 0x1340
		x"60",x"67",x"67",x"00",x"FF",x"63",x"28",x"30", -- 0x1348
		x"0E",x"0C",x"15",x"76",x"0F",x"4C",x"6C",x"2E", -- 0x1350
		x"E7",x"F1",x"FF",x"FF",x"7F",x"BF",x"DF",x"E0", -- 0x1358
		x"31",x"8F",x"E7",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x1360
		x"63",x"45",x"20",x"E8",x"76",x"18",x"C7",x"FF", -- 0x1368
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"14",x"F8", -- 0x1370
		x"B0",x"14",x"0B",x"A4",x"CF",x"66",x"11",x"FF", -- 0x1378
		x"FF",x"F9",x"F0",x"E8",x"D1",x"D4",x"E8",x"B5", -- 0x1380
		x"9F",x"D9",x"C8",x"E8",x"E5",x"E6",x"E9",x"F3", -- 0x1388
		x"FF",x"FF",x"AC",x"40",x"49",x"A4",x"C0",x"F6", -- 0x1390
		x"BE",x"9E",x"FF",x"3F",x"3F",x"38",x"BF",x"BF", -- 0x1398
		x"C9",x"E9",x"E4",x"F3",x"FF",x"FF",x"FF",x"EF", -- 0x13A0
		x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF", -- 0x13A8
		x"BF",x"BF",x"BF",x"C1",x"FE",x"FE",x"FE",x"FE", -- 0x13B0
		x"FE",x"1F",x"E7",x"F3",x"A3",x"41",x"51",x"20", -- 0x13B8
		x"EF",x"EE",x"EE",x"EF",x"EF",x"EF",x"EF",x"EF", -- 0x13C0
		x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF", -- 0x13C8
		x"EA",x"D2",x"42",x"66",x"6E",x"3E",x"BE",x"9E", -- 0x13D0
		x"FF",x"C0",x"DF",x"DC",x"DF",x"DF",x"DF",x"DF", -- 0x13D8
		x"F8",x"E8",x"E4",x"FA",x"E4",x"F8",x"D9",x"D6", -- 0x13E0
		x"D5",x"CE",x"EA",x"E7",x"F2",x"FB",x"FF",x"FF", -- 0x13E8
		x"5D",x"DD",x"5C",x"5E",x"1E",x"1F",x"1F",x"5F", -- 0x13F0
		x"5E",x"41",x"87",x"D0",x"6A",x"1D",x"C3",x"FF", -- 0x13F8
		x"AA",x"5B",x"56",x"BB",x"AC",x"56",x"EA",x"FF", -- 0x1400
		x"D5",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1408
		x"AA",x"34",x"52",x"34",x"55",x"88",x"DE",x"F5", -- 0x1410
		x"7F",x"56",x"80",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1418
		x"4B",x"EA",x"5B",x"74",x"C9",x"69",x"32",x"B3", -- 0x1420
		x"EA",x"D5",x"FF",x"D5",x"FF",x"FF",x"FF",x"FF", -- 0x1428
		x"AA",x"BB",x"56",x"94",x"2F",x"94",x"BA",x"55", -- 0x1430
		x"AD",x"5D",x"EA",x"7F",x"E5",x"FF",x"FF",x"FF", -- 0x1438
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1440
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1448
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1450
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1458
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1460
		x"FF",x"FF",x"FF",x"FF",x"FC",x"FA",x"F9",x"FB", -- 0x1468
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1470
		x"FF",x"FF",x"FF",x"FF",x"7F",x"E3",x"47",x"27", -- 0x1478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"81", -- 0x1480
		x"BC",x"46",x"E3",x"07",x"24",x"25",x"9D",x"D4", -- 0x1488
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"81", -- 0x1490
		x"01",x"46",x"3A",x"2A",x"42",x"22",x"5B",x"7B", -- 0x1498
		x"00",x"01",x"AA",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x14A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14A8
		x"00",x"55",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14B8
		x"AA",x"A5",x"94",x"56",x"34",x"49",x"2E",x"13", -- 0x14C0
		x"95",x"8D",x"43",x"20",x"90",x"C9",x"E8",x"E4", -- 0x14C8
		x"AA",x"71",x"1A",x"DD",x"29",x"D2",x"FC",x"2B", -- 0x14D0
		x"55",x"6E",x"15",x"79",x"CE",x"4D",x"54",x"25", -- 0x14D8
		x"FA",x"FD",x"FD",x"FE",x"FE",x"FF",x"FF",x"CF", -- 0x14E0
		x"CF",x"FF",x"83",x"FF",x"E7",x"E7",x"E7",x"E7", -- 0x14E8
		x"2E",x"35",x"16",x"8F",x"9B",x"44",x"8A",x"A3", -- 0x14F0
		x"D7",x"D0",x"D3",x"E9",x"E8",x"F5",x"F4",x"F4", -- 0x14F8
		x"55",x"93",x"6C",x"95",x"2F",x"D9",x"AA",x"FF", -- 0x1500
		x"D7",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1508
		x"55",x"AA",x"AD",x"0B",x"50",x"5A",x"D2",x"FF", -- 0x1510
		x"2A",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1518
		x"55",x"AA",x"2A",x"54",x"9A",x"6B",x"35",x"AD", -- 0x1520
		x"A4",x"FF",x"55",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1528
		x"55",x"BB",x"0A",x"56",x"A5",x"A9",x"7A",x"96", -- 0x1530
		x"AA",x"FF",x"55",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1538
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1540
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1548
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1550
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1558
		x"AA",x"54",x"51",x"A8",x"00",x"55",x"00",x"FF", -- 0x1560
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1568
		x"B4",x"AA",x"49",x"54",x"43",x"00",x"55",x"00", -- 0x1570
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1578
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1580
		x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x1588
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1590
		x"FF",x"80",x"3E",x"42",x"2A",x"82",x"2A",x"5A", -- 0x1598
		x"FE",x"00",x"AA",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x15A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15A8
		x"00",x"00",x"AA",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x15B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E8
		x"9C",x"9C",x"9C",x"9C",x"9C",x"9C",x"9C",x"9C", -- 0x15F0
		x"9C",x"9F",x"9F",x"9F",x"9F",x"FF",x"FF",x"FF", -- 0x15F8
		x"55",x"AA",x"D9",x"D5",x"FF",x"FF",x"FF",x"00", -- 0x1600
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1608
		x"54",x"BB",x"A9",x"56",x"DA",x"D1",x"FF",x"7F", -- 0x1610
		x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1618
		x"55",x"EB",x"4A",x"2D",x"98",x"A6",x"55",x"AA", -- 0x1620
		x"EA",x"BF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1628
		x"55",x"AA",x"CA",x"3B",x"D4",x"49",x"B6",x"A4", -- 0x1630
		x"AB",x"FF",x"D5",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1640
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FA",x"F5", -- 0x1648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1650
		x"FE",x"FD",x"F6",x"C9",x"37",x"E8",x"D6",x"59", -- 0x1658
		x"99",x"1B",x"08",x"CC",x"E6",x"00",x"FF",x"FF", -- 0x1660
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1668
		x"14",x"1A",x"85",x"E4",x"77",x"21",x"80",x"FF", -- 0x1670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1680
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1688
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1690
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1698
		x"55",x"A2",x"00",x"AA",x"00",x"FF",x"FF",x"FF", -- 0x16A0
		x"FF",x"FF",x"FF",x"FF",x"FC",x"FA",x"F9",x"FB", -- 0x16A8
		x"FF",x"80",x"2A",x"80",x"7F",x"FF",x"FF",x"FF", -- 0x16B0
		x"FF",x"FF",x"FF",x"FF",x"7F",x"E3",x"47",x"27", -- 0x16B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16D8
		x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x16E0
		x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x16E8
		x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07", -- 0x16F0
		x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07", -- 0x16F8
		x"55",x"AB",x"1A",x"66",x"7F",x"FF",x"F5",x"C0", -- 0x1700
		x"FF",x"DF",x"FF",x"DF",x"FF",x"DF",x"FF",x"DF", -- 0x1708
		x"55",x"4A",x"93",x"36",x"FF",x"FF",x"55",x"00", -- 0x1710
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1718
		x"45",x"B4",x"CA",x"B5",x"57",x"6E",x"5B",x"A4", -- 0x1720
		x"FF",x"55",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1728
		x"55",x"AA",x"CB",x"65",x"5A",x"A9",x"AA",x"92", -- 0x1730
		x"FF",x"55",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1738
		x"55",x"EC",x"4A",x"D5",x"49",x"2A",x"22",x"BA", -- 0x1740
		x"55",x"FF",x"8A",x"FF",x"BE",x"FF",x"FF",x"FF", -- 0x1748
		x"55",x"EE",x"91",x"62",x"5C",x"A9",x"D4",x"15", -- 0x1750
		x"6C",x"A2",x"CD",x"56",x"FF",x"5B",x"FF",x"FF", -- 0x1758
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1760
		x"FF",x"FF",x"FF",x"FF",x"FF",x"C7",x"AE",x"84", -- 0x1768
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"7F", -- 0x1778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1788
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1790
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1798
		x"55",x"AB",x"65",x"D8",x"01",x"56",x"01",x"FF", -- 0x17A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"C7",x"AE",x"84", -- 0x17A8
		x"55",x"2A",x"BB",x"00",x"55",x"00",x"FF",x"FF", -- 0x17B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"7F", -- 0x17B8
		x"4A",x"95",x"A0",x"64",x"41",x"D5",x"AA",x"2B", -- 0x17C0
		x"DE",x"28",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x17C8
		x"8A",x"55",x"25",x"8B",x"59",x"2B",x"DB",x"67", -- 0x17D0
		x"87",x"07",x"07",x"07",x"07",x"07",x"07",x"07", -- 0x17D8
		x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",x"FE",x"FF", -- 0x17E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E8
		x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"87", -- 0x17F0
		x"E7",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1800
		x"FF",x"FF",x"FF",x"00",x"AA",x"00",x"FF",x"FF", -- 0x1808
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1810
		x"FF",x"FF",x"FF",x"7F",x"80",x"2A",x"80",x"9C", -- 0x1818
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1820
		x"FF",x"00",x"56",x"01",x"FC",x"FF",x"FF",x"FF", -- 0x1828
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1830
		x"FF",x"FF",x"00",x"55",x"00",x"FF",x"FF",x"FF", -- 0x1838
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1840
		x"FF",x"00",x"55",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1848
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1850
		x"00",x"55",x"00",x"3F",x"FF",x"FF",x"FF",x"FF", -- 0x1858
		x"7F",x"5F",x"7F",x"5F",x"7F",x"5F",x"7F",x"1F", -- 0x1860
		x"00",x"3B",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1868
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1870
		x"00",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1878
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1880
		x"EF",x"EF",x"EF",x"EF",x"E7",x"03",x"FF",x"FF", -- 0x1888
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1890
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1898
		x"2F",x"EF",x"FF",x"AF",x"AF",x"AF",x"CF",x"9F", -- 0x18A0
		x"2F",x"4F",x"C0",x"F7",x"F5",x"F6",x"63",x"8F", -- 0x18A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18B0
		x"FF",x"80",x"39",x"7F",x"FF",x"F7",x"1F",x"FF", -- 0x18B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18D8
		x"FE",x"02",x"C2",x"82",x"82",x"CA",x"7A",x"B0", -- 0x18E0
		x"C1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18E8
		x"FE",x"02",x"22",x"A2",x"A2",x"9A",x"82",x"F9", -- 0x18F0
		x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18F8
		x"AA",x"54",x"51",x"A8",x"2A",x"D4",x"AC",x"2A", -- 0x1900
		x"D4",x"AA",x"00",x"54",x"01",x"F8",x"FF",x"FF", -- 0x1908
		x"B4",x"AA",x"49",x"54",x"83",x"88",x"44",x"55", -- 0x1910
		x"9A",x"82",x"21",x"05",x"50",x"05",x"E0",x"FF", -- 0x1918
		x"FF",x"FF",x"FF",x"07",x"03",x"F1",x"F8",x"FC", -- 0x1920
		x"3E",x"1F",x"8F",x"C7",x"E7",x"E7",x"E7",x"E7", -- 0x1928
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x1930
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x1938
		x"C7",x"C7",x"C7",x"E7",x"C7",x"8F",x"1F",x"3E", -- 0x1940
		x"FC",x"F8",x"F1",x"03",x"07",x"FF",x"FF",x"FF", -- 0x1948
		x"17",x"17",x"17",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x1950
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1958
		x"FF",x"FF",x"F8",x"01",x"54",x"00",x"FC",x"F9", -- 0x1960
		x"F9",x"F2",x"F4",x"E9",x"E2",x"C9",x"E5",x"14", -- 0x1968
		x"FF",x"E0",x"05",x"50",x"03",x"84",x"B2",x"4D", -- 0x1970
		x"68",x"4A",x"95",x"52",x"54",x"29",x"4A",x"B4", -- 0x1978
		x"FF",x"FF",x"FF",x"9F",x"47",x"C7",x"80",x"FF", -- 0x1980
		x"FF",x"1F",x"DD",x"DF",x"EB",x"E8",x"EB",x"6A", -- 0x1988
		x"FF",x"FF",x"FF",x"CF",x"A3",x"E1",x"C1",x"FE", -- 0x1990
		x"FE",x"1E",x"86",x"F2",x"FE",x"0E",x"E7",x"EF", -- 0x1998
		x"28",x"2B",x"AB",x"29",x"2C",x"6E",x"EF",x"EF", -- 0x19A0
		x"CF",x"9B",x"33",x"70",x"67",x"FE",x"00",x"00", -- 0x19A8
		x"00",x"C1",x"63",x"9C",x"FA",x"05",x"FD",x"FE", -- 0x19B0
		x"F5",x"E8",x"D0",x"27",x"4F",x"9C",x"38",x"70", -- 0x19B8
		x"03",x"FE",x"01",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19C8
		x"E6",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19D8
		x"FE",x"FC",x"FC",x"FD",x"FD",x"FC",x"FE",x"FF", -- 0x19E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19E8
		x"FE",x"AA",x"AA",x"6A",x"6E",x"BE",x"60",x"01", -- 0x19F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19F8
		x"AA",x"54",x"51",x"A8",x"2A",x"D4",x"2A",x"FF", -- 0x1A00
		x"80",x"2A",x"80",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A08
		x"B4",x"AA",x"49",x"54",x"83",x"88",x"44",x"55", -- 0x1A10
		x"FF",x"00",x"2A",x"80",x"FF",x"FF",x"FF",x"FF", -- 0x1A18
		x"FF",x"FF",x"FF",x"0F",x"07",x"E3",x"F0",x"F8", -- 0x1A20
		x"3C",x"1F",x"8F",x"C7",x"E7",x"E7",x"E7",x"E7", -- 0x1A28
		x"FF",x"FF",x"FF",x"C0",x"80",x"1F",x"3F",x"7F", -- 0x1A30
		x"F0",x"E0",x"C7",x"8F",x"9F",x"9F",x"9F",x"9F", -- 0x1A38
		x"C7",x"C7",x"C7",x"E7",x"C7",x"8F",x"1F",x"3C", -- 0x1A40
		x"F8",x"F0",x"E3",x"07",x"0F",x"FF",x"FF",x"FF", -- 0x1A48
		x"8F",x"8F",x"8F",x"9F",x"8F",x"C7",x"E0",x"F0", -- 0x1A50
		x"7F",x"3F",x"1F",x"80",x"C0",x"FF",x"FF",x"FF", -- 0x1A58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"2A",x"80", -- 0x1A60
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A68
		x"FF",x"FF",x"FF",x"FF",x"80",x"2A",x"00",x"FF", -- 0x1A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A78
		x"8F",x"C7",x"03",x"FF",x"FF",x"FF",x"FC",x"FF", -- 0x1A80
		x"A7",x"BF",x"BF",x"89",x"87",x"87",x"AE",x"AE", -- 0x1A88
		x"FF",x"FF",x"FF",x"FF",x"80",x"FF",x"00",x"FF", -- 0x1A90
		x"03",x"FE",x"FF",x"FF",x"FF",x"FE",x"7E",x"F7", -- 0x1A98
		x"AE",x"AE",x"AE",x"A6",x"A6",x"B3",x"B8",x"BC", -- 0x1AA0
		x"23",x"19",x"00",x"00",x"0F",x"07",x"80",x"00", -- 0x1AA8
		x"A7",x"C7",x"AB",x"73",x"03",x"FE",x"F8",x"03", -- 0x1AB0
		x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00", -- 0x1AB8
		x"20",x"00",x"9F",x"00",x"3F",x"FF",x"FF",x"FF", -- 0x1AC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AC8
		x"00",x"00",x"00",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x1AD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AD8
		x"F8",x"F5",x"F0",x"F4",x"FE",x"FD",x"FC",x"F8", -- 0x1AE0
		x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AE8
		x"FF",x"C7",x"8F",x"4F",x"5F",x"2F",x"0F",x"5F", -- 0x1AF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AF8
		x"AA",x"54",x"51",x"A8",x"2A",x"03",x"50",x"05", -- 0x1B00
		x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B08
		x"B4",x"AA",x"49",x"54",x"83",x"55",x"4B",x"00", -- 0x1B10
		x"55",x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8", -- 0x1B20
		x"F1",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3",x"F3", -- 0x1B28
		x"FF",x"FF",x"FF",x"80",x"00",x"3F",x"7F",x"FF", -- 0x1B30
		x"F0",x"E0",x"C7",x"8F",x"9F",x"9F",x"9F",x"9F", -- 0x1B38
		x"E3",x"E3",x"E3",x"F3",x"F3",x"F3",x"F3",x"F1", -- 0x1B40
		x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B48
		x"8F",x"8F",x"8F",x"9F",x"8F",x"C7",x"E0",x"F0", -- 0x1B50
		x"FF",x"7F",x"3F",x"00",x"80",x"FF",x"FF",x"FF", -- 0x1B58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0", -- 0x1B60
		x"05",x"50",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"55", -- 0x1B70
		x"00",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B78
		x"FF",x"00",x"00",x"80",x"70",x"1C",x"04",x"C0", -- 0x1B80
		x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B88
		x"FF",x"00",x"00",x"00",x"0B",x"CF",x"CF",x"CE", -- 0x1B90
		x"CF",x"40",x"1C",x"22",x"3D",x"9E",x"17",x"17", -- 0x1B98
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"0C", -- 0x1BA0
		x"F0",x"00",x"EB",x"19",x"04",x"06",x"23",x"93", -- 0x1BA8
		x"57",x"57",x"57",x"D1",x"87",x"17",x"17",x"16", -- 0x1BB0
		x"97",x"57",x"17",x"C5",x"90",x"05",x"02",x"06", -- 0x1BB8
		x"78",x"3C",x"1F",x"0F",x"00",x"FF",x"FF",x"FF", -- 0x1BC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BC8
		x"00",x"03",x"FF",x"FF",x"00",x"FF",x"FF",x"FF", -- 0x1BD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"5F",x"2F",x"AB", -- 0x1BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x1FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
