-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_M6 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_M6 is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"60",x"80",x"0A",x"81",x"C4",x"81",x"7E",x"82", -- 0x0000
		x"1C",x"83",x"D8",x"83",x"94",x"84",x"61",x"85", -- 0x0008
		x"FD",x"85",x"B7",x"86",x"77",x"87",x"69",x"88", -- 0x0010
		x"19",x"89",x"D5",x"89",x"B3",x"8A",x"C8",x"8B", -- 0x0018
		x"68",x"8C",x"24",x"8D",x"F8",x"8D",x"EA",x"8E", -- 0x0020
		x"88",x"8F",x"9E",x"90",x"A8",x"91",x"D1",x"92", -- 0x0028
		x"73",x"93",x"61",x"94",x"75",x"95",x"8D",x"96", -- 0x0030
		x"2F",x"97",x"31",x"98",x"37",x"99",x"70",x"9A", -- 0x0038
		x"68",x"8C",x"24",x"8D",x"F8",x"8D",x"EA",x"8E", -- 0x0040
		x"88",x"8F",x"9E",x"90",x"A8",x"91",x"D1",x"92", -- 0x0048
		x"73",x"93",x"61",x"94",x"75",x"95",x"8D",x"96", -- 0x0050
		x"2F",x"97",x"31",x"98",x"37",x"99",x"70",x"9A", -- 0x0058
		x"80",x"C0",x"FE",x"FE",x"FD",x"84",x"C1",x"20", -- 0x0060
		x"00",x"FE",x"20",x"00",x"FE",x"FD",x"84",x"C2", -- 0x0068
		x"20",x"00",x"03",x"11",x"FE",x"20",x"00",x"FE", -- 0x0070
		x"FD",x"84",x"C3",x"20",x"00",x"FE",x"20",x"00", -- 0x0078
		x"FE",x"FD",x"84",x"C2",x"00",x"03",x"00",x"04", -- 0x0080
		x"10",x"21",x"FE",x"00",x"03",x"00",x"04",x"FE", -- 0x0088
		x"FD",x"84",x"C2",x"00",x"03",x"00",x"04",x"FE", -- 0x0090
		x"00",x"03",x"00",x"04",x"08",x"00",x"FE",x"FD", -- 0x0098
		x"84",x"C2",x"00",x"03",x"00",x"04",x"FE",x"00", -- 0x00A0
		x"03",x"00",x"04",x"FE",x"FD",x"85",x"C2",x"00", -- 0x00A8
		x"03",x"00",x"04",x"FE",x"03",x"11",x"00",x"03", -- 0x00B0
		x"00",x"04",x"FE",x"FD",x"85",x"C2",x"00",x"03", -- 0x00B8
		x"00",x"04",x"FE",x"00",x"03",x"00",x"04",x"FE", -- 0x00C0
		x"FD",x"85",x"C3",x"00",x"03",x"00",x"04",x"10", -- 0x00C8
		x"21",x"FE",x"03",x"11",x"00",x"03",x"00",x"04", -- 0x00D0
		x"FE",x"FD",x"85",x"C3",x"00",x"03",x"00",x"04", -- 0x00D8
		x"FE",x"00",x"03",x"00",x"04",x"FE",x"FD",x"84", -- 0x00E0
		x"C3",x"08",x"00",x"20",x"00",x"FE",x"20",x"00", -- 0x00E8
		x"FE",x"FD",x"84",x"C3",x"20",x"01",x"20",x"02", -- 0x00F0
		x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD",x"83", -- 0x00F8
		x"C0",x"20",x"01",x"20",x"02",x"FE",x"FE",x"FD", -- 0x0100
		x"FC",x"FF",x"80",x"C0",x"FE",x"FE",x"FD",x"84", -- 0x0108
		x"C2",x"20",x"01",x"20",x"02",x"FE",x"20",x"01", -- 0x0110
		x"20",x"02",x"FE",x"FD",x"84",x"C2",x"20",x"01", -- 0x0118
		x"20",x"02",x"23",x"11",x"FE",x"20",x"01",x"20", -- 0x0120
		x"02",x"FE",x"FD",x"84",x"C3",x"20",x"01",x"20", -- 0x0128
		x"02",x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x0130
		x"84",x"C3",x"20",x"01",x"20",x"02",x"10",x"20", -- 0x0138
		x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD",x"84", -- 0x0140
		x"C3",x"00",x"10",x"00",x"11",x"FE",x"08",x"00", -- 0x0148
		x"00",x"10",x"00",x"11",x"FE",x"FD",x"84",x"C3", -- 0x0150
		x"00",x"10",x"00",x"11",x"FE",x"00",x"10",x"00", -- 0x0158
		x"11",x"FE",x"FD",x"84",x"C3",x"00",x"10",x"00", -- 0x0160
		x"11",x"23",x"11",x"FE",x"00",x"10",x"00",x"11", -- 0x0168
		x"FE",x"FD",x"85",x"C3",x"00",x"10",x"00",x"11", -- 0x0170
		x"FE",x"00",x"10",x"00",x"11",x"FE",x"FD",x"85", -- 0x0178
		x"C3",x"00",x"03",x"00",x"04",x"10",x"20",x"FE", -- 0x0180
		x"00",x"03",x"00",x"04",x"03",x"12",x"FE",x"FD", -- 0x0188
		x"85",x"C3",x"00",x"03",x"00",x"04",x"FE",x"00", -- 0x0190
		x"03",x"00",x"04",x"FE",x"FD",x"84",x"C3",x"08", -- 0x0198
		x"00",x"20",x"01",x"20",x"02",x"FE",x"20",x"01", -- 0x01A0
		x"20",x"02",x"FE",x"FD",x"84",x"C3",x"20",x"01", -- 0x01A8
		x"20",x"02",x"FE",x"20",x"01",x"20",x"02",x"FE", -- 0x01B0
		x"FD",x"83",x"C0",x"20",x"01",x"20",x"02",x"FE", -- 0x01B8
		x"FE",x"FD",x"FC",x"FF",x"80",x"C0",x"FE",x"FE", -- 0x01C0
		x"FD",x"84",x"C3",x"20",x"1A",x"20",x"1B",x"FE", -- 0x01C8
		x"20",x"1A",x"20",x"1B",x"FE",x"FD",x"84",x"C3", -- 0x01D0
		x"20",x"1A",x"20",x"1B",x"03",x"12",x"FE",x"20", -- 0x01D8
		x"1A",x"20",x"1B",x"FE",x"FD",x"84",x"C3",x"20", -- 0x01E0
		x"1A",x"20",x"1B",x"FE",x"20",x"1A",x"20",x"1B", -- 0x01E8
		x"FE",x"FD",x"84",x"C3",x"00",x"12",x"00",x"13", -- 0x01F0
		x"10",x"22",x"FE",x"00",x"12",x"00",x"13",x"FE", -- 0x01F8
		x"FD",x"85",x"C3",x"00",x"12",x"00",x"13",x"FE", -- 0x0200
		x"08",x"00",x"00",x"12",x"00",x"13",x"FE",x"FD", -- 0x0208
		x"85",x"C3",x"00",x"12",x"00",x"13",x"FE",x"00", -- 0x0210
		x"12",x"00",x"13",x"FE",x"FD",x"85",x"C3",x"00", -- 0x0218
		x"12",x"00",x"13",x"23",x"12",x"FE",x"00",x"12", -- 0x0220
		x"00",x"13",x"FE",x"FD",x"85",x"C4",x"00",x"12", -- 0x0228
		x"00",x"13",x"FE",x"00",x"12",x"00",x"13",x"FE", -- 0x0230
		x"FD",x"85",x"C4",x"00",x"12",x"00",x"13",x"10", -- 0x0238
		x"22",x"FE",x"23",x"12",x"00",x"12",x"00",x"13", -- 0x0240
		x"FE",x"FD",x"85",x"C4",x"00",x"12",x"00",x"13", -- 0x0248
		x"FE",x"00",x"03",x"00",x"04",x"FE",x"FD",x"85", -- 0x0250
		x"C4",x"08",x"00",x"20",x"01",x"20",x"02",x"FE", -- 0x0258
		x"20",x"01",x"20",x"02",x"FE",x"FD",x"85",x"C3", -- 0x0260
		x"20",x"01",x"20",x"02",x"FE",x"20",x"01",x"20", -- 0x0268
		x"02",x"FE",x"FD",x"84",x"C0",x"20",x"01",x"20", -- 0x0270
		x"02",x"FE",x"FE",x"FD",x"FC",x"FF",x"80",x"C0", -- 0x0278
		x"FE",x"FE",x"FD",x"85",x"C0",x"20",x"00",x"FE", -- 0x0280
		x"20",x"00",x"FE",x"FD",x"85",x"C0",x"20",x"00", -- 0x0288
		x"FE",x"20",x"00",x"FE",x"FD",x"85",x"C0",x"20", -- 0x0290
		x"00",x"FE",x"20",x"00",x"FE",x"FD",x"85",x"C0", -- 0x0298
		x"20",x"00",x"FE",x"03",x"A0",x"FE",x"FD",x"85", -- 0x02A0
		x"C0",x"20",x"01",x"20",x"02",x"FE",x"20",x"01", -- 0x02A8
		x"20",x"02",x"FE",x"FD",x"86",x"C0",x"20",x"01", -- 0x02B0
		x"20",x"02",x"FE",x"20",x"01",x"20",x"02",x"10", -- 0x02B8
		x"61",x"FE",x"FD",x"86",x"C0",x"20",x"01",x"20", -- 0x02C0
		x"02",x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x02C8
		x"86",x"C0",x"20",x"01",x"20",x"02",x"FE",x"03", -- 0x02D0
		x"C1",x"FE",x"FD",x"86",x"C0",x"20",x"1A",x"20", -- 0x02D8
		x"1B",x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD", -- 0x02E0
		x"86",x"C0",x"20",x"1A",x"20",x"1B",x"FE",x"20", -- 0x02E8
		x"1A",x"20",x"1B",x"FE",x"FD",x"85",x"C0",x"08", -- 0x02F0
		x"00",x"20",x"1A",x"20",x"1B",x"FE",x"20",x"1A", -- 0x02F8
		x"20",x"1B",x"FE",x"FD",x"85",x"C0",x"20",x"1A", -- 0x0300
		x"20",x"1B",x"FE",x"20",x"1A",x"20",x"1B",x"FE", -- 0x0308
		x"FD",x"83",x"C0",x"20",x"1A",x"20",x"1B",x"FE", -- 0x0310
		x"FE",x"FD",x"FC",x"FF",x"80",x"C0",x"FE",x"FE", -- 0x0318
		x"FD",x"85",x"C3",x"20",x"1C",x"20",x"1D",x"FE", -- 0x0320
		x"20",x"1C",x"20",x"1D",x"FE",x"FD",x"85",x"C3", -- 0x0328
		x"20",x"1C",x"20",x"1D",x"03",x"12",x"FE",x"20", -- 0x0330
		x"1C",x"20",x"1D",x"FE",x"FD",x"86",x"C3",x"20", -- 0x0338
		x"1C",x"20",x"1D",x"FE",x"20",x"1C",x"20",x"1D", -- 0x0340
		x"FE",x"FD",x"86",x"C3",x"20",x"1C",x"20",x"1D", -- 0x0348
		x"10",x"21",x"FE",x"20",x"1C",x"20",x"1D",x"FE", -- 0x0350
		x"FD",x"86",x"C4",x"00",x"14",x"00",x"15",x"08", -- 0x0358
		x"00",x"FE",x"00",x"14",x"00",x"15",x"FE",x"FD", -- 0x0360
		x"86",x"C4",x"00",x"14",x"00",x"15",x"FE",x"00", -- 0x0368
		x"14",x"00",x"15",x"FE",x"FD",x"86",x"C4",x"00", -- 0x0370
		x"14",x"00",x"15",x"03",x"82",x"FE",x"00",x"14", -- 0x0378
		x"00",x"15",x"FE",x"FD",x"86",x"C4",x"00",x"14", -- 0x0380
		x"00",x"15",x"FE",x"00",x"14",x"00",x"15",x"FE", -- 0x0388
		x"FD",x"86",x"C5",x"00",x"14",x"00",x"15",x"10", -- 0x0390
		x"21",x"FE",x"00",x"14",x"00",x"15",x"03",x"A3", -- 0x0398
		x"FE",x"FD",x"87",x"C5",x"02",x"00",x"20",x"00", -- 0x03A0
		x"FE",x"02",x"00",x"20",x"00",x"FE",x"FD",x"86", -- 0x03A8
		x"C4",x"08",x"00",x"02",x"00",x"FE",x"20",x"00", -- 0x03B0
		x"20",x"00",x"02",x"00",x"20",x"00",x"FE",x"FD", -- 0x03B8
		x"85",x"C4",x"02",x"00",x"20",x"00",x"FE",x"02", -- 0x03C0
		x"00",x"20",x"00",x"FE",x"FD",x"84",x"C0",x"02", -- 0x03C8
		x"00",x"20",x"00",x"FE",x"FE",x"FD",x"FC",x"FF", -- 0x03D0
		x"80",x"C0",x"FE",x"FE",x"FD",x"86",x"C4",x"20", -- 0x03D8
		x"00",x"FE",x"20",x"00",x"10",x"24",x"FE",x"FD", -- 0x03E0
		x"86",x"C4",x"20",x"00",x"03",x"AC",x"FE",x"20", -- 0x03E8
		x"00",x"FE",x"FD",x"86",x"C4",x"00",x"16",x"00", -- 0x03F0
		x"17",x"FE",x"00",x"16",x"00",x"17",x"FE",x"FD", -- 0x03F8
		x"86",x"C4",x"00",x"16",x"00",x"17",x"10",x"23", -- 0x0400
		x"FE",x"00",x"16",x"00",x"17",x"FE",x"FD",x"86", -- 0x0408
		x"C5",x"00",x"16",x"00",x"17",x"FE",x"00",x"16", -- 0x0410
		x"00",x"17",x"08",x"00",x"FE",x"FD",x"86",x"C5", -- 0x0418
		x"00",x"16",x"00",x"17",x"FE",x"00",x"16",x"00", -- 0x0420
		x"17",x"FE",x"FD",x"86",x"C5",x"00",x"16",x"00", -- 0x0428
		x"17",x"20",x"00",x"03",x"CD",x"FE",x"00",x"16", -- 0x0430
		x"00",x"17",x"20",x"00",x"FE",x"FD",x"86",x"C5", -- 0x0438
		x"00",x"16",x"00",x"17",x"20",x"00",x"FE",x"00", -- 0x0440
		x"16",x"00",x"17",x"20",x"00",x"FE",x"FD",x"87", -- 0x0448
		x"C5",x"00",x"16",x"00",x"17",x"10",x"23",x"FE", -- 0x0450
		x"00",x"16",x"00",x"17",x"03",x"CE",x"FE",x"FD", -- 0x0458
		x"86",x"C4",x"01",x"03",x"01",x"04",x"FE",x"01", -- 0x0460
		x"03",x"01",x"04",x"FE",x"FD",x"86",x"C3",x"01", -- 0x0468
		x"03",x"01",x"04",x"08",x"00",x"FE",x"01",x"03", -- 0x0470
		x"01",x"04",x"FE",x"FD",x"85",x"C3",x"01",x"03", -- 0x0478
		x"01",x"04",x"FE",x"01",x"03",x"01",x"04",x"FE", -- 0x0480
		x"FD",x"84",x"C0",x"01",x"03",x"01",x"04",x"FE", -- 0x0488
		x"FE",x"FD",x"FC",x"FF",x"80",x"C0",x"FE",x"FE", -- 0x0490
		x"FD",x"86",x"C4",x"20",x"1D",x"20",x"1E",x"FE", -- 0x0498
		x"20",x"1D",x"20",x"1E",x"FE",x"FD",x"86",x"C4", -- 0x04A0
		x"20",x"1D",x"20",x"1E",x"23",x"C7",x"FE",x"20", -- 0x04A8
		x"1D",x"20",x"1E",x"FE",x"FD",x"86",x"C4",x"20", -- 0x04B0
		x"1D",x"20",x"1E",x"FE",x"20",x"1D",x"20",x"1E", -- 0x04B8
		x"FE",x"FD",x"86",x"C4",x"00",x"14",x"00",x"15", -- 0x04C0
		x"10",x"22",x"FE",x"00",x"14",x"00",x"15",x"FE", -- 0x04C8
		x"FD",x"86",x"C5",x"00",x"14",x"00",x"15",x"08", -- 0x04D0
		x"00",x"FE",x"00",x"14",x"00",x"15",x"FE",x"FD", -- 0x04D8
		x"86",x"C5",x"00",x"14",x"00",x"15",x"FE",x"00", -- 0x04E0
		x"14",x"00",x"15",x"FE",x"FD",x"86",x"C5",x"00", -- 0x04E8
		x"14",x"00",x"15",x"20",x"01",x"20",x"02",x"23", -- 0x04F0
		x"C8",x"FE",x"00",x"14",x"00",x"15",x"20",x"01", -- 0x04F8
		x"20",x"02",x"FE",x"FD",x"86",x"C5",x"00",x"14", -- 0x0500
		x"00",x"15",x"20",x"01",x"20",x"02",x"FE",x"00", -- 0x0508
		x"14",x"00",x"15",x"20",x"01",x"20",x"02",x"FE", -- 0x0510
		x"FD",x"87",x"C5",x"00",x"14",x"00",x"15",x"10", -- 0x0518
		x"22",x"FE",x"00",x"14",x"00",x"15",x"23",x"C1", -- 0x0520
		x"FE",x"FD",x"87",x"C5",x"00",x"03",x"00",x"04", -- 0x0528
		x"FE",x"00",x"03",x"00",x"04",x"FE",x"FD",x"86", -- 0x0530
		x"C4",x"00",x"03",x"00",x"04",x"28",x"00",x"FE", -- 0x0538
		x"00",x"03",x"00",x"04",x"FE",x"FD",x"85",x"C4", -- 0x0540
		x"00",x"03",x"00",x"04",x"FE",x"00",x"03",x"00", -- 0x0548
		x"04",x"FE",x"FD",x"84",x"C0",x"00",x"03",x"00", -- 0x0550
		x"04",x"FE",x"FE",x"FD",x"09",x"00",x"FD",x"FC", -- 0x0558
		x"FF",x"80",x"C0",x"FE",x"FE",x"FD",x"85",x"C0", -- 0x0560
		x"20",x"1A",x"20",x"1B",x"FE",x"20",x"1A",x"20", -- 0x0568
		x"1B",x"FE",x"FD",x"85",x"C0",x"20",x"1A",x"20", -- 0x0570
		x"1B",x"10",x"63",x"FE",x"20",x"1A",x"20",x"1B", -- 0x0578
		x"FE",x"FD",x"85",x"C0",x"20",x"1A",x"20",x"1B", -- 0x0580
		x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD",x"85", -- 0x0588
		x"C0",x"20",x"1A",x"20",x"1B",x"FE",x"23",x"C2", -- 0x0590
		x"FE",x"FD",x"86",x"C0",x"20",x"1C",x"20",x"1D", -- 0x0598
		x"FE",x"20",x"1C",x"20",x"1D",x"FE",x"FD",x"86", -- 0x05A0
		x"C0",x"20",x"1C",x"20",x"1D",x"10",x"66",x"FE", -- 0x05A8
		x"20",x"1C",x"20",x"1D",x"FE",x"FD",x"87",x"C0", -- 0x05B0
		x"20",x"1C",x"20",x"1D",x"FE",x"20",x"1C",x"20", -- 0x05B8
		x"1D",x"FE",x"FD",x"87",x"C0",x"20",x"1C",x"20", -- 0x05C0
		x"1D",x"FE",x"03",x"EB",x"FE",x"FD",x"87",x"C0", -- 0x05C8
		x"20",x"00",x"FE",x"20",x"00",x"FE",x"FD",x"86", -- 0x05D0
		x"C0",x"20",x"00",x"FE",x"20",x"00",x"FE",x"FD", -- 0x05D8
		x"85",x"C0",x"28",x"00",x"20",x"00",x"FE",x"20", -- 0x05E0
		x"00",x"FE",x"FD",x"85",x"C0",x"20",x"00",x"FE", -- 0x05E8
		x"20",x"00",x"FE",x"FD",x"83",x"C0",x"20",x"00", -- 0x05F0
		x"FE",x"FE",x"FD",x"FC",x"FF",x"80",x"C0",x"FE", -- 0x05F8
		x"FE",x"FD",x"84",x"D2",x"20",x"1A",x"20",x"1B", -- 0x0600
		x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD",x"84", -- 0x0608
		x"D2",x"20",x"1A",x"20",x"1B",x"03",x"A4",x"FE", -- 0x0610
		x"20",x"1A",x"20",x"1B",x"FE",x"FD",x"85",x"D2", -- 0x0618
		x"20",x"1A",x"20",x"1B",x"FE",x"20",x"1A",x"20", -- 0x0620
		x"1B",x"FE",x"FD",x"85",x"D2",x"10",x"21",x"20", -- 0x0628
		x"1A",x"20",x"1B",x"FE",x"20",x"1A",x"20",x"1B", -- 0x0630
		x"FE",x"FD",x"85",x"D2",x"00",x"12",x"00",x"13", -- 0x0638
		x"FE",x"00",x"12",x"00",x"13",x"08",x"00",x"FE", -- 0x0640
		x"FD",x"85",x"D3",x"00",x"12",x"00",x"13",x"FE", -- 0x0648
		x"00",x"12",x"00",x"13",x"FE",x"FD",x"85",x"D3", -- 0x0650
		x"00",x"12",x"00",x"13",x"03",x"CD",x"FE",x"00", -- 0x0658
		x"12",x"00",x"13",x"FE",x"FD",x"86",x"D3",x"00", -- 0x0660
		x"12",x"00",x"13",x"FE",x"00",x"12",x"00",x"13", -- 0x0668
		x"FE",x"FD",x"86",x"D3",x"00",x"12",x"00",x"13", -- 0x0670
		x"10",x"21",x"FE",x"00",x"12",x"00",x"13",x"03", -- 0x0678
		x"D6",x"FE",x"FD",x"87",x"D3",x"20",x"1E",x"20", -- 0x0680
		x"1F",x"FE",x"20",x"1E",x"20",x"1F",x"FE",x"FD", -- 0x0688
		x"86",x"D2",x"20",x"1E",x"20",x"1F",x"08",x"00", -- 0x0690
		x"FE",x"20",x"1E",x"20",x"1F",x"FE",x"FD",x"85", -- 0x0698
		x"D2",x"20",x"1E",x"20",x"1F",x"FE",x"20",x"1E", -- 0x06A0
		x"20",x"1F",x"FE",x"FD",x"84",x"D0",x"20",x"1E", -- 0x06A8
		x"20",x"1F",x"FE",x"FE",x"FD",x"FC",x"FF",x"80", -- 0x06B0
		x"C0",x"FE",x"FE",x"FD",x"85",x"D3",x"20",x"00", -- 0x06B8
		x"FE",x"20",x"00",x"FE",x"FD",x"85",x"D4",x"20", -- 0x06C0
		x"00",x"FE",x"03",x"CF",x"20",x"00",x"FE",x"FD", -- 0x06C8
		x"86",x"D4",x"20",x"01",x"20",x"02",x"FE",x"20", -- 0x06D0
		x"01",x"20",x"02",x"FE",x"FD",x"86",x"D4",x"20", -- 0x06D8
		x"01",x"20",x"02",x"10",x"65",x"FE",x"20",x"01", -- 0x06E0
		x"20",x"02",x"FE",x"FD",x"86",x"D4",x"20",x"18", -- 0x06E8
		x"20",x"19",x"FE",x"08",x"00",x"20",x"18",x"20", -- 0x06F0
		x"19",x"FE",x"FD",x"86",x"D4",x"01",x"03",x"01", -- 0x06F8
		x"04",x"FE",x"01",x"03",x"01",x"04",x"FE",x"FD", -- 0x0700
		x"86",x"D5",x"01",x"03",x"01",x"04",x"FE",x"23", -- 0x0708
		x"C0",x"01",x"03",x"01",x"04",x"FE",x"FD",x"86", -- 0x0710
		x"D5",x"01",x"03",x"01",x"04",x"FE",x"01",x"03", -- 0x0718
		x"01",x"04",x"FE",x"FD",x"86",x"D5",x"10",x"65", -- 0x0720
		x"01",x"03",x"01",x"04",x"FE",x"23",x"E1",x"01", -- 0x0728
		x"03",x"01",x"04",x"FE",x"FD",x"87",x"D5",x"22", -- 0x0730
		x"00",x"00",x"12",x"00",x"13",x"FE",x"22",x"00", -- 0x0738
		x"00",x"12",x"00",x"13",x"FE",x"FD",x"86",x"D4", -- 0x0740
		x"22",x"00",x"28",x"00",x"00",x"12",x"00",x"13", -- 0x0748
		x"FE",x"22",x"00",x"00",x"12",x"00",x"13",x"FE", -- 0x0750
		x"FD",x"85",x"D4",x"00",x"12",x"00",x"13",x"22", -- 0x0758
		x"00",x"FE",x"00",x"12",x"00",x"13",x"22",x"00", -- 0x0760
		x"FE",x"FD",x"84",x"D0",x"00",x"12",x"00",x"13", -- 0x0768
		x"22",x"00",x"FE",x"FE",x"FD",x"FC",x"FF",x"80", -- 0x0770
		x"C0",x"FE",x"FE",x"FD",x"85",x"D4",x"20",x"1A", -- 0x0778
		x"20",x"1B",x"FE",x"20",x"1A",x"20",x"1B",x"FE", -- 0x0780
		x"FD",x"85",x"D4",x"20",x"1A",x"20",x"1B",x"23", -- 0x0788
		x"CB",x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD", -- 0x0790
		x"85",x"D4",x"20",x"1A",x"20",x"1B",x"FE",x"20", -- 0x0798
		x"1A",x"20",x"1B",x"FE",x"FD",x"86",x"D4",x"20", -- 0x07A0
		x"1A",x"20",x"1B",x"10",x"22",x"FE",x"20",x"1A", -- 0x07A8
		x"20",x"1B",x"FE",x"FD",x"86",x"D4",x"00",x"10", -- 0x07B0
		x"00",x"11",x"21",x"12",x"21",x"13",x"28",x"00", -- 0x07B8
		x"FE",x"00",x"10",x"00",x"11",x"21",x"12",x"21", -- 0x07C0
		x"13",x"FE",x"FD",x"86",x"D4",x"00",x"10",x"00", -- 0x07C8
		x"11",x"21",x"12",x"21",x"13",x"FE",x"00",x"10", -- 0x07D0
		x"00",x"11",x"21",x"12",x"21",x"13",x"FE",x"FD", -- 0x07D8
		x"86",x"D5",x"00",x"10",x"00",x"11",x"21",x"12", -- 0x07E0
		x"21",x"13",x"23",x"D4",x"FE",x"00",x"10",x"00", -- 0x07E8
		x"11",x"21",x"12",x"21",x"13",x"FE",x"FD",x"86", -- 0x07F0
		x"D5",x"01",x"12",x"01",x"13",x"20",x"1C",x"20", -- 0x07F8
		x"1D",x"FE",x"20",x"1C",x"20",x"1D",x"01",x"12", -- 0x0800
		x"01",x"13",x"FE",x"FD",x"87",x"D5",x"20",x"1C", -- 0x0808
		x"20",x"1D",x"01",x"12",x"01",x"13",x"10",x"22", -- 0x0810
		x"FE",x"20",x"1C",x"20",x"1D",x"01",x"12",x"01", -- 0x0818
		x"13",x"23",x"EC",x"FE",x"FD",x"87",x"D5",x"04", -- 0x0820
		x"03",x"20",x"1C",x"20",x"1D",x"FE",x"20",x"1C", -- 0x0828
		x"20",x"1D",x"04",x"40",x"FE",x"FD",x"86",x"D4", -- 0x0830
		x"04",x"03",x"20",x"1C",x"20",x"1D",x"FE",x"20", -- 0x0838
		x"1C",x"20",x"1D",x"28",x"00",x"04",x"40",x"FE", -- 0x0840
		x"FD",x"86",x"D3",x"04",x"03",x"20",x"1C",x"20", -- 0x0848
		x"1D",x"FE",x"20",x"1C",x"20",x"1D",x"FE",x"04", -- 0x0850
		x"40",x"FD",x"85",x"D2",x"04",x"03",x"20",x"1C", -- 0x0858
		x"20",x"1D",x"FE",x"FE",x"04",x"40",x"FD",x"FC", -- 0x0860
		x"FF",x"80",x"C0",x"FE",x"FE",x"FD",x"85",x"C0", -- 0x0868
		x"20",x"01",x"20",x"02",x"FE",x"20",x"01",x"20", -- 0x0870
		x"02",x"FE",x"FD",x"85",x"C0",x"20",x"01",x"20", -- 0x0878
		x"02",x"10",x"67",x"FE",x"20",x"01",x"20",x"02", -- 0x0880
		x"FE",x"FD",x"85",x"C0",x"20",x"01",x"20",x"02", -- 0x0888
		x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD",x"85", -- 0x0890
		x"C0",x"20",x"01",x"20",x"02",x"FE",x"23",x"CD", -- 0x0898
		x"FE",x"FD",x"85",x"C0",x"20",x"01",x"20",x"02", -- 0x08A0
		x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD",x"85", -- 0x08A8
		x"C0",x"20",x"01",x"20",x"02",x"10",x"64",x"FE", -- 0x08B0
		x"20",x"01",x"20",x"02",x"FE",x"FD",x"85",x"C0", -- 0x08B8
		x"20",x"01",x"20",x"02",x"FE",x"20",x"01",x"20", -- 0x08C0
		x"02",x"FE",x"FD",x"86",x"C0",x"20",x"01",x"20", -- 0x08C8
		x"02",x"FE",x"23",x"E6",x"FE",x"FD",x"86",x"C0", -- 0x08D0
		x"20",x"01",x"20",x"02",x"FE",x"20",x"01",x"20", -- 0x08D8
		x"02",x"FE",x"FD",x"86",x"C0",x"20",x"01",x"20", -- 0x08E0
		x"02",x"10",x"20",x"FE",x"20",x"01",x"20",x"02", -- 0x08E8
		x"FE",x"FD",x"84",x"C0",x"20",x"01",x"20",x"02", -- 0x08F0
		x"28",x"00",x"FE",x"20",x"01",x"20",x"02",x"FE", -- 0x08F8
		x"FD",x"85",x"C0",x"20",x"01",x"20",x"02",x"FE", -- 0x0900
		x"20",x"01",x"20",x"02",x"FE",x"FD",x"83",x"C0", -- 0x0908
		x"20",x"01",x"20",x"02",x"FE",x"FE",x"FD",x"FC", -- 0x0910
		x"FF",x"80",x"C0",x"FE",x"FE",x"FD",x"86",x"D3", -- 0x0918
		x"20",x"1C",x"20",x"1D",x"FE",x"20",x"1C",x"20", -- 0x0920
		x"1D",x"10",x"24",x"FE",x"FD",x"86",x"D3",x"20", -- 0x0928
		x"1C",x"20",x"1D",x"23",x"B0",x"FE",x"20",x"1C", -- 0x0930
		x"20",x"1D",x"FE",x"FD",x"86",x"D4",x"20",x"1C", -- 0x0938
		x"20",x"1D",x"FE",x"20",x"1C",x"20",x"1D",x"FE", -- 0x0940
		x"FD",x"86",x"D4",x"00",x"12",x"00",x"13",x"10", -- 0x0948
		x"21",x"FE",x"00",x"12",x"00",x"13",x"FE",x"FD", -- 0x0950
		x"86",x"D4",x"00",x"12",x"00",x"13",x"28",x"00", -- 0x0958
		x"FE",x"00",x"12",x"00",x"13",x"FE",x"FD",x"86", -- 0x0960
		x"D4",x"00",x"12",x"00",x"13",x"FE",x"00",x"12", -- 0x0968
		x"00",x"13",x"FE",x"FD",x"86",x"D4",x"00",x"12", -- 0x0970
		x"00",x"13",x"23",x"C9",x"FE",x"00",x"12",x"00", -- 0x0978
		x"13",x"FE",x"FD",x"87",x"D4",x"20",x"18",x"20", -- 0x0980
		x"19",x"FE",x"20",x"18",x"20",x"19",x"FE",x"FD", -- 0x0988
		x"87",x"D4",x"20",x"18",x"20",x"19",x"10",x"21", -- 0x0990
		x"FE",x"03",x"D2",x"20",x"18",x"20",x"19",x"FE", -- 0x0998
		x"FD",x"87",x"D4",x"20",x"18",x"20",x"19",x"FE", -- 0x09A0
		x"20",x"18",x"20",x"19",x"FE",x"FD",x"87",x"D4", -- 0x09A8
		x"20",x"18",x"20",x"19",x"28",x"00",x"FE",x"20", -- 0x09B0
		x"18",x"20",x"19",x"FE",x"FD",x"85",x"D4",x"20", -- 0x09B8
		x"18",x"20",x"19",x"FE",x"20",x"18",x"20",x"19", -- 0x09C0
		x"FE",x"FD",x"84",x"D2",x"20",x"18",x"20",x"19", -- 0x09C8
		x"FE",x"FE",x"FD",x"FC",x"FF",x"80",x"C0",x"FE", -- 0x09D0
		x"FE",x"FD",x"87",x"D3",x"01",x"03",x"01",x"04", -- 0x09D8
		x"FE",x"01",x"03",x"01",x"04",x"FE",x"FD",x"87", -- 0x09E0
		x"D3",x"01",x"03",x"01",x"04",x"23",x"CB",x"FE", -- 0x09E8
		x"01",x"03",x"01",x"04",x"FE",x"FD",x"87",x"D3", -- 0x09F0
		x"01",x"03",x"01",x"04",x"FE",x"20",x"1A",x"20", -- 0x09F8
		x"1B",x"FE",x"FD",x"87",x"D4",x"20",x"1A",x"20", -- 0x0A00
		x"1B",x"10",x"20",x"FE",x"20",x"1A",x"20",x"1B", -- 0x0A08
		x"FE",x"FD",x"87",x"D4",x"20",x"1A",x"20",x"1B", -- 0x0A10
		x"28",x"00",x"FE",x"20",x"1A",x"20",x"1B",x"FE", -- 0x0A18
		x"FD",x"87",x"D4",x"20",x"1A",x"20",x"1B",x"FE", -- 0x0A20
		x"00",x"12",x"00",x"13",x"FE",x"FD",x"87",x"D4", -- 0x0A28
		x"00",x"12",x"00",x"13",x"23",x"CC",x"FE",x"00", -- 0x0A30
		x"12",x"00",x"13",x"FE",x"FD",x"88",x"D4",x"00", -- 0x0A38
		x"12",x"00",x"13",x"FE",x"00",x"12",x"00",x"13", -- 0x0A40
		x"FE",x"FD",x"88",x"D4",x"00",x"16",x"00",x"17", -- 0x0A48
		x"20",x"01",x"20",x"02",x"10",x"20",x"FE",x"00", -- 0x0A50
		x"16",x"00",x"17",x"20",x"01",x"20",x"02",x"23", -- 0x0A58
		x"E5",x"FE",x"FD",x"88",x"D4",x"00",x"16",x"00", -- 0x0A60
		x"17",x"20",x"01",x"20",x"02",x"FE",x"00",x"16", -- 0x0A68
		x"00",x"17",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x0A70
		x"88",x"D4",x"00",x"16",x"00",x"17",x"20",x"01", -- 0x0A78
		x"20",x"02",x"28",x"00",x"FE",x"00",x"16",x"00", -- 0x0A80
		x"17",x"20",x"01",x"20",x"02",x"FE",x"FD",x"86", -- 0x0A88
		x"D4",x"00",x"16",x"00",x"17",x"20",x"01",x"20", -- 0x0A90
		x"02",x"FE",x"00",x"16",x"00",x"17",x"20",x"01", -- 0x0A98
		x"20",x"02",x"FE",x"FD",x"85",x"D3",x"00",x"16", -- 0x0AA0
		x"00",x"17",x"20",x"01",x"20",x"02",x"FE",x"FE", -- 0x0AA8
		x"FD",x"FC",x"FF",x"80",x"C0",x"FE",x"FE",x"FD", -- 0x0AB0
		x"87",x"E4",x"00",x"16",x"00",x"17",x"20",x"00", -- 0x0AB8
		x"FE",x"00",x"16",x"00",x"17",x"20",x"00",x"FE", -- 0x0AC0
		x"FD",x"87",x"E4",x"00",x"16",x"00",x"17",x"20", -- 0x0AC8
		x"00",x"23",x"E6",x"FE",x"00",x"16",x"00",x"17", -- 0x0AD0
		x"20",x"00",x"FE",x"FD",x"87",x"E4",x"00",x"16", -- 0x0AD8
		x"00",x"17",x"20",x"00",x"FE",x"00",x"16",x"00", -- 0x0AE0
		x"17",x"20",x"00",x"FE",x"FD",x"88",x"E4",x"00", -- 0x0AE8
		x"16",x"00",x"17",x"20",x"01",x"20",x"02",x"10", -- 0x0AF0
		x"65",x"FE",x"00",x"16",x"00",x"17",x"20",x"01", -- 0x0AF8
		x"20",x"02",x"FE",x"FD",x"88",x"E4",x"00",x"16", -- 0x0B00
		x"00",x"17",x"20",x"01",x"20",x"02",x"28",x"00", -- 0x0B08
		x"FE",x"00",x"16",x"00",x"17",x"20",x"01",x"20", -- 0x0B10
		x"02",x"FE",x"FD",x"88",x"E4",x"00",x"16",x"00", -- 0x0B18
		x"17",x"20",x"01",x"20",x"02",x"FE",x"00",x"16", -- 0x0B20
		x"00",x"17",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x0B28
		x"88",x"E4",x"00",x"16",x"00",x"17",x"20",x"01", -- 0x0B30
		x"20",x"02",x"23",x"E8",x"FE",x"00",x"16",x"00", -- 0x0B38
		x"17",x"20",x"01",x"20",x"02",x"FE",x"FD",x"88", -- 0x0B40
		x"E4",x"00",x"10",x"00",x"11",x"20",x"1C",x"20", -- 0x0B48
		x"1D",x"FE",x"00",x"10",x"00",x"11",x"20",x"1C", -- 0x0B50
		x"20",x"1D",x"FE",x"FD",x"88",x"E5",x"00",x"10", -- 0x0B58
		x"00",x"11",x"20",x"1C",x"20",x"1D",x"10",x"20", -- 0x0B60
		x"FE",x"23",x"F0",x"00",x"10",x"00",x"11",x"20", -- 0x0B68
		x"1C",x"20",x"1D",x"FE",x"FD",x"88",x"E5",x"00", -- 0x0B70
		x"10",x"00",x"11",x"20",x"1C",x"20",x"1D",x"FE", -- 0x0B78
		x"00",x"10",x"00",x"11",x"20",x"1C",x"20",x"1D", -- 0x0B80
		x"FE",x"FD",x"88",x"E5",x"00",x"10",x"00",x"11", -- 0x0B88
		x"20",x"1E",x"20",x"1F",x"28",x"00",x"FE",x"00", -- 0x0B90
		x"10",x"00",x"11",x"20",x"1E",x"20",x"1F",x"FE", -- 0x0B98
		x"FD",x"86",x"E4",x"00",x"10",x"00",x"11",x"20", -- 0x0BA0
		x"1E",x"20",x"1F",x"FE",x"00",x"10",x"00",x"11", -- 0x0BA8
		x"20",x"1E",x"20",x"1F",x"FE",x"FD",x"85",x"E3", -- 0x0BB0
		x"00",x"10",x"00",x"11",x"20",x"1E",x"20",x"1F", -- 0x0BB8
		x"FE",x"FE",x"FD",x"09",x"00",x"FD",x"FC",x"FF", -- 0x0BC0
		x"80",x"C0",x"FE",x"FE",x"FD",x"85",x"C0",x"10", -- 0x0BC8
		x"60",x"FE",x"10",x"61",x"FE",x"FD",x"85",x"C0", -- 0x0BD0
		x"23",x"E9",x"FE",x"FE",x"FD",x"85",x"C0",x"20", -- 0x0BD8
		x"00",x"FE",x"20",x"00",x"FE",x"FD",x"85",x"C0", -- 0x0BE0
		x"20",x"00",x"28",x"00",x"FE",x"20",x"00",x"FE", -- 0x0BE8
		x"FD",x"85",x"C0",x"20",x"00",x"FE",x"20",x"00", -- 0x0BF0
		x"FE",x"FD",x"85",x"C0",x"20",x"01",x"20",x"02", -- 0x0BF8
		x"10",x"62",x"FE",x"20",x"01",x"20",x"02",x"10", -- 0x0C00
		x"65",x"FE",x"FD",x"85",x"C0",x"10",x"63",x"20", -- 0x0C08
		x"01",x"20",x"02",x"FE",x"20",x"01",x"20",x"02", -- 0x0C10
		x"FE",x"FD",x"85",x"C0",x"20",x"01",x"20",x"02", -- 0x0C18
		x"23",x"F2",x"FE",x"20",x"01",x"20",x"02",x"FE", -- 0x0C20
		x"FD",x"86",x"C0",x"20",x"01",x"20",x"02",x"FE", -- 0x0C28
		x"10",x"65",x"FE",x"FD",x"86",x"C0",x"20",x"1A", -- 0x0C30
		x"20",x"1B",x"FE",x"20",x"1A",x"20",x"1B",x"FE", -- 0x0C38
		x"FD",x"85",x"C0",x"20",x"1A",x"20",x"1B",x"28", -- 0x0C40
		x"00",x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD", -- 0x0C48
		x"85",x"C0",x"20",x"1A",x"20",x"1B",x"FE",x"20", -- 0x0C50
		x"1A",x"20",x"1B",x"FE",x"FD",x"83",x"C0",x"20", -- 0x0C58
		x"1A",x"20",x"1B",x"FE",x"FE",x"FD",x"FC",x"FF", -- 0x0C60
		x"80",x"C0",x"FE",x"FE",x"FD",x"85",x"D2",x"00", -- 0x0C68
		x"14",x"00",x"15",x"FE",x"00",x"14",x"00",x"15", -- 0x0C70
		x"FE",x"FD",x"85",x"D2",x"00",x"14",x"00",x"15", -- 0x0C78
		x"23",x"12",x"FE",x"00",x"14",x"00",x"15",x"FE", -- 0x0C80
		x"FD",x"85",x"D2",x"00",x"14",x"00",x"15",x"FE", -- 0x0C88
		x"00",x"14",x"00",x"15",x"FE",x"FD",x"85",x"D2", -- 0x0C90
		x"00",x"14",x"00",x"15",x"10",x"21",x"FE",x"00", -- 0x0C98
		x"14",x"00",x"15",x"FE",x"FD",x"85",x"D2",x"00", -- 0x0CA0
		x"14",x"00",x"15",x"28",x"00",x"FE",x"00",x"14", -- 0x0CA8
		x"00",x"15",x"FE",x"FD",x"85",x"D3",x"00",x"14", -- 0x0CB0
		x"00",x"15",x"FE",x"00",x"14",x"00",x"15",x"FE", -- 0x0CB8
		x"FD",x"85",x"D3",x"00",x"14",x"00",x"15",x"23", -- 0x0CC0
		x"12",x"FE",x"00",x"14",x"00",x"15",x"FE",x"FD", -- 0x0CC8
		x"85",x"D3",x"20",x"1B",x"04",x"04",x"FE",x"20", -- 0x0CD0
		x"1B",x"04",x"40",x"FE",x"FD",x"86",x"D3",x"20", -- 0x0CD8
		x"1B",x"10",x"21",x"04",x"04",x"FE",x"23",x"D3", -- 0x0CE0
		x"20",x"1B",x"04",x"40",x"FE",x"FD",x"86",x"D3", -- 0x0CE8
		x"20",x"1B",x"04",x"04",x"FE",x"20",x"1B",x"04", -- 0x0CF0
		x"40",x"FE",x"FD",x"84",x"D2",x"20",x"1B",x"28", -- 0x0CF8
		x"00",x"04",x"04",x"FE",x"20",x"1B",x"04",x"40", -- 0x0D00
		x"FE",x"FD",x"85",x"D2",x"20",x"1B",x"04",x"04", -- 0x0D08
		x"FE",x"20",x"1B",x"04",x"40",x"FE",x"FD",x"84", -- 0x0D10
		x"D0",x"20",x"1B",x"04",x"04",x"FE",x"04",x"40", -- 0x0D18
		x"FE",x"FD",x"FC",x"FF",x"80",x"C0",x"FE",x"FE", -- 0x0D20
		x"FD",x"86",x"D3",x"04",x"03",x"FE",x"04",x"40", -- 0x0D28
		x"10",x"24",x"FE",x"FD",x"86",x"D3",x"03",x"B4", -- 0x0D30
		x"04",x"03",x"FE",x"20",x"00",x"04",x"40",x"FE", -- 0x0D38
		x"FD",x"86",x"D4",x"04",x"03",x"20",x"00",x"FE", -- 0x0D40
		x"20",x"00",x"04",x"40",x"FE",x"FD",x"86",x"D4", -- 0x0D48
		x"10",x"23",x"04",x"03",x"20",x"00",x"FE",x"20", -- 0x0D50
		x"00",x"04",x"40",x"FE",x"FD",x"86",x"D4",x"28", -- 0x0D58
		x"00",x"04",x"04",x"20",x"01",x"20",x"02",x"FE", -- 0x0D60
		x"20",x"01",x"20",x"02",x"04",x"40",x"FE",x"FD", -- 0x0D68
		x"86",x"D4",x"04",x"04",x"20",x"01",x"20",x"02", -- 0x0D70
		x"FE",x"20",x"01",x"20",x"02",x"04",x"40",x"FE", -- 0x0D78
		x"FD",x"86",x"D4",x"23",x"CD",x"04",x"04",x"20", -- 0x0D80
		x"01",x"20",x"02",x"FE",x"20",x"01",x"20",x"02", -- 0x0D88
		x"04",x"40",x"FE",x"FD",x"86",x"D4",x"04",x"04", -- 0x0D90
		x"20",x"01",x"20",x"02",x"FE",x"20",x"01",x"20", -- 0x0D98
		x"02",x"04",x"40",x"FE",x"FD",x"86",x"D4",x"10", -- 0x0DA0
		x"23",x"22",x"01",x"04",x"04",x"FE",x"23",x"D6", -- 0x0DA8
		x"22",x"01",x"04",x"40",x"FE",x"FD",x"86",x"D4", -- 0x0DB0
		x"22",x"01",x"04",x"04",x"20",x"00",x"FE",x"22", -- 0x0DB8
		x"01",x"20",x"00",x"04",x"40",x"FE",x"FD",x"86", -- 0x0DC0
		x"D4",x"22",x"01",x"28",x"00",x"04",x"04",x"FE", -- 0x0DC8
		x"22",x"01",x"20",x"00",x"04",x"40",x"FE",x"FD", -- 0x0DD0
		x"86",x"D3",x"22",x"01",x"04",x"04",x"20",x"00", -- 0x0DD8
		x"FE",x"22",x"01",x"20",x"00",x"04",x"40",x"FE", -- 0x0DE0
		x"FD",x"84",x"D0",x"22",x"01",x"04",x"04",x"20", -- 0x0DE8
		x"00",x"FE",x"FE",x"04",x"40",x"FD",x"FC",x"FF", -- 0x0DF0
		x"80",x"C0",x"FE",x"FE",x"FD",x"86",x"D3",x"20", -- 0x0DF8
		x"18",x"20",x"19",x"FE",x"20",x"18",x"20",x"19", -- 0x0E00
		x"FE",x"FD",x"86",x"D3",x"23",x"C7",x"20",x"18", -- 0x0E08
		x"20",x"19",x"FE",x"20",x"18",x"20",x"19",x"FE", -- 0x0E10
		x"FD",x"86",x"D4",x"20",x"18",x"20",x"19",x"FE", -- 0x0E18
		x"20",x"18",x"20",x"19",x"FE",x"FD",x"86",x"D4", -- 0x0E20
		x"20",x"18",x"20",x"19",x"10",x"22",x"FE",x"20", -- 0x0E28
		x"18",x"20",x"19",x"FE",x"FD",x"86",x"D5",x"20", -- 0x0E30
		x"18",x"20",x"19",x"28",x"00",x"FE",x"20",x"18", -- 0x0E38
		x"20",x"19",x"FE",x"FD",x"86",x"D5",x"20",x"18", -- 0x0E40
		x"20",x"19",x"20",x"01",x"20",x"02",x"FE",x"20", -- 0x0E48
		x"18",x"20",x"19",x"20",x"01",x"20",x"02",x"FE", -- 0x0E50
		x"FD",x"86",x"D6",x"20",x"18",x"20",x"19",x"20", -- 0x0E58
		x"01",x"20",x"02",x"23",x"C8",x"FE",x"20",x"18", -- 0x0E60
		x"20",x"19",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x0E68
		x"86",x"D6",x"00",x"16",x"00",x"17",x"20",x"01", -- 0x0E70
		x"20",x"02",x"FE",x"00",x"16",x"00",x"17",x"20", -- 0x0E78
		x"01",x"20",x"02",x"FE",x"FD",x"86",x"D6",x"00", -- 0x0E80
		x"16",x"00",x"17",x"20",x"1A",x"20",x"1B",x"10", -- 0x0E88
		x"22",x"FE",x"23",x"D1",x"00",x"16",x"00",x"17", -- 0x0E90
		x"20",x"1A",x"20",x"1B",x"FE",x"FD",x"86",x"D6", -- 0x0E98
		x"00",x"16",x"00",x"17",x"20",x"1A",x"20",x"1B", -- 0x0EA0
		x"FE",x"00",x"16",x"00",x"17",x"20",x"1A",x"20", -- 0x0EA8
		x"1B",x"FE",x"FD",x"86",x"D5",x"28",x"00",x"00", -- 0x0EB0
		x"16",x"00",x"17",x"20",x"1A",x"20",x"1B",x"FE", -- 0x0EB8
		x"00",x"16",x"00",x"17",x"20",x"1A",x"20",x"1B", -- 0x0EC0
		x"FE",x"FD",x"87",x"D6",x"00",x"16",x"00",x"17", -- 0x0EC8
		x"20",x"1A",x"20",x"1B",x"FE",x"00",x"16",x"00", -- 0x0ED0
		x"17",x"20",x"00",x"FE",x"FD",x"86",x"D0",x"00", -- 0x0ED8
		x"16",x"00",x"17",x"20",x"00",x"FE",x"FE",x"FD", -- 0x0EE0
		x"FC",x"FF",x"80",x"C0",x"FE",x"FE",x"FD",x"85", -- 0x0EE8
		x"C0",x"23",x"E2",x"FE",x"20",x"00",x"FE",x"FD", -- 0x0EF0
		x"85",x"C0",x"20",x"00",x"FE",x"20",x"00",x"FE", -- 0x0EF8
		x"FD",x"85",x"C0",x"20",x"00",x"10",x"66",x"FE", -- 0x0F00
		x"20",x"00",x"FE",x"FD",x"85",x"C0",x"20",x"00", -- 0x0F08
		x"10",x"63",x"FE",x"20",x"00",x"FE",x"FD",x"86", -- 0x0F10
		x"C0",x"10",x"65",x"FE",x"10",x"62",x"FE",x"FD", -- 0x0F18
		x"86",x"C0",x"20",x"01",x"20",x"02",x"FE",x"20", -- 0x0F20
		x"01",x"20",x"02",x"FE",x"FD",x"86",x"C0",x"20", -- 0x0F28
		x"01",x"20",x"02",x"FE",x"20",x"01",x"20",x"02", -- 0x0F30
		x"23",x"C9",x"FE",x"FD",x"86",x"C0",x"20",x"01", -- 0x0F38
		x"20",x"02",x"FE",x"20",x"01",x"20",x"02",x"FE", -- 0x0F40
		x"FD",x"86",x"C0",x"23",x"D3",x"FE",x"20",x"1A", -- 0x0F48
		x"20",x"1B",x"FE",x"FD",x"86",x"C0",x"20",x"1A", -- 0x0F50
		x"20",x"1B",x"FE",x"20",x"1A",x"20",x"1B",x"FE", -- 0x0F58
		x"FD",x"85",x"C0",x"20",x"1A",x"20",x"1B",x"28", -- 0x0F60
		x"00",x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD", -- 0x0F68
		x"85",x"C0",x"20",x"1A",x"20",x"1B",x"FE",x"20", -- 0x0F70
		x"1A",x"20",x"1B",x"FE",x"FD",x"84",x"C0",x"20", -- 0x0F78
		x"1A",x"20",x"1B",x"FE",x"FE",x"FD",x"FC",x"FF", -- 0x0F80
		x"80",x"C4",x"FE",x"FE",x"FD",x"84",x"D2",x"00", -- 0x0F88
		x"10",x"00",x"11",x"20",x"01",x"20",x"02",x"FE", -- 0x0F90
		x"00",x"10",x"00",x"11",x"20",x"01",x"20",x"02", -- 0x0F98
		x"FE",x"FD",x"84",x"D2",x"00",x"10",x"00",x"11", -- 0x0FA0
		x"20",x"01",x"20",x"02",x"23",x"12",x"FE",x"00", -- 0x0FA8
		x"10",x"00",x"11",x"20",x"01",x"20",x"02",x"FE", -- 0x0FB0
		x"FD",x"84",x"D3",x"00",x"10",x"00",x"11",x"20", -- 0x0FB8
		x"01",x"20",x"02",x"FE",x"00",x"10",x"00",x"11", -- 0x0FC0
		x"20",x"01",x"20",x"02",x"FE",x"FD",x"84",x"D3", -- 0x0FC8
		x"00",x"10",x"00",x"11",x"20",x"01",x"20",x"02", -- 0x0FD0
		x"10",x"21",x"FE",x"00",x"10",x"00",x"11",x"20", -- 0x0FD8
		x"01",x"20",x"02",x"FE",x"FD",x"85",x"D3",x"00", -- 0x0FE0
		x"10",x"00",x"11",x"20",x"01",x"20",x"02",x"28", -- 0x0FE8
		x"00",x"FE",x"00",x"10",x"00",x"11",x"20",x"01", -- 0x0FF0
		x"20",x"02",x"FE",x"FD",x"85",x"D3",x"00",x"10", -- 0x0FF8
		x"00",x"11",x"20",x"01",x"20",x"02",x"FE",x"00", -- 0x1000
		x"10",x"00",x"11",x"20",x"01",x"20",x"02",x"FE", -- 0x1008
		x"FD",x"85",x"D3",x"00",x"10",x"00",x"11",x"20", -- 0x1010
		x"01",x"20",x"02",x"23",x"CC",x"FE",x"00",x"10", -- 0x1018
		x"00",x"11",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x1020
		x"85",x"D3",x"01",x"12",x"01",x"13",x"20",x"1C", -- 0x1028
		x"20",x"1D",x"FE",x"01",x"12",x"01",x"13",x"20", -- 0x1030
		x"1C",x"20",x"1D",x"FE",x"FD",x"85",x"D3",x"01", -- 0x1038
		x"12",x"01",x"13",x"20",x"1C",x"20",x"1D",x"10", -- 0x1040
		x"21",x"FE",x"23",x"D5",x"01",x"12",x"01",x"13", -- 0x1048
		x"20",x"1C",x"20",x"1D",x"FE",x"FD",x"85",x"D3", -- 0x1050
		x"01",x"12",x"01",x"13",x"20",x"1C",x"20",x"1D", -- 0x1058
		x"FE",x"01",x"12",x"01",x"13",x"20",x"1C",x"20", -- 0x1060
		x"1D",x"FE",x"FD",x"85",x"D3",x"01",x"12",x"01", -- 0x1068
		x"13",x"20",x"1C",x"20",x"1D",x"28",x"00",x"FE", -- 0x1070
		x"01",x"12",x"01",x"13",x"20",x"1C",x"20",x"1D", -- 0x1078
		x"FE",x"FD",x"85",x"D3",x"01",x"12",x"01",x"13", -- 0x1080
		x"20",x"1C",x"20",x"1D",x"FE",x"01",x"12",x"01", -- 0x1088
		x"13",x"FE",x"FD",x"84",x"D2",x"01",x"12",x"01", -- 0x1090
		x"13",x"FE",x"FE",x"FD",x"FC",x"FF",x"80",x"C0", -- 0x1098
		x"FE",x"FE",x"FD",x"86",x"D3",x"21",x"03",x"21", -- 0x10A0
		x"04",x"FE",x"21",x"03",x"21",x"04",x"FE",x"FD", -- 0x10A8
		x"86",x"D3",x"21",x"03",x"21",x"04",x"FE",x"21", -- 0x10B0
		x"03",x"21",x"04",x"03",x"D6",x"FE",x"FD",x"86", -- 0x10B8
		x"D3",x"21",x"03",x"21",x"04",x"20",x"01",x"20", -- 0x10C0
		x"02",x"FE",x"21",x"03",x"21",x"04",x"20",x"01", -- 0x10C8
		x"20",x"02",x"FE",x"FD",x"86",x"D4",x"21",x"03", -- 0x10D0
		x"21",x"04",x"20",x"01",x"20",x"02",x"FE",x"21", -- 0x10D8
		x"03",x"21",x"04",x"20",x"01",x"20",x"02",x"10", -- 0x10E0
		x"20",x"FE",x"FD",x"86",x"D4",x"00",x"12",x"00", -- 0x10E8
		x"13",x"20",x"01",x"20",x"02",x"28",x"00",x"FE", -- 0x10F0
		x"00",x"12",x"00",x"13",x"20",x"01",x"20",x"02", -- 0x10F8
		x"FE",x"FD",x"86",x"D4",x"00",x"12",x"00",x"13", -- 0x1100
		x"20",x"01",x"20",x"02",x"FE",x"00",x"12",x"00", -- 0x1108
		x"13",x"20",x"01",x"20",x"02",x"FE",x"FD",x"86", -- 0x1110
		x"D5",x"00",x"12",x"00",x"13",x"20",x"01",x"20", -- 0x1118
		x"02",x"23",x"E7",x"FE",x"00",x"12",x"00",x"13", -- 0x1120
		x"20",x"01",x"20",x"02",x"FE",x"FD",x"86",x"D5", -- 0x1128
		x"00",x"12",x"00",x"13",x"20",x"01",x"20",x"02", -- 0x1130
		x"FE",x"00",x"12",x"00",x"13",x"20",x"01",x"20", -- 0x1138
		x"02",x"FE",x"FD",x"87",x"D5",x"20",x"1C",x"20", -- 0x1140
		x"1D",x"00",x"10",x"00",x"11",x"10",x"20",x"FE", -- 0x1148
		x"03",x"E8",x"20",x"1C",x"20",x"1D",x"00",x"10", -- 0x1150
		x"00",x"11",x"FE",x"FD",x"87",x"D5",x"20",x"1C", -- 0x1158
		x"20",x"1D",x"00",x"10",x"00",x"11",x"FE",x"20", -- 0x1160
		x"1C",x"20",x"1D",x"00",x"10",x"00",x"11",x"FE", -- 0x1168
		x"FD",x"87",x"D5",x"20",x"1C",x"20",x"1D",x"22", -- 0x1170
		x"01",x"28",x"00",x"FE",x"20",x"1C",x"20",x"1D", -- 0x1178
		x"22",x"01",x"FE",x"FD",x"86",x"D4",x"20",x"1C", -- 0x1180
		x"20",x"1D",x"00",x"10",x"00",x"11",x"FE",x"20", -- 0x1188
		x"1C",x"20",x"1D",x"00",x"10",x"00",x"11",x"FE", -- 0x1190
		x"FD",x"85",x"D3",x"20",x"1C",x"20",x"1D",x"00", -- 0x1198
		x"10",x"00",x"11",x"FE",x"FE",x"FD",x"FC",x"FF", -- 0x11A0
		x"80",x"C0",x"FE",x"FE",x"FD",x"87",x"E4",x"20", -- 0x11A8
		x"00",x"01",x"14",x"01",x"15",x"FE",x"20",x"00", -- 0x11B0
		x"01",x"14",x"01",x"15",x"FE",x"FD",x"87",x"E4", -- 0x11B8
		x"20",x"00",x"01",x"14",x"01",x"15",x"23",x"E1", -- 0x11C0
		x"FE",x"20",x"00",x"01",x"14",x"01",x"15",x"FE", -- 0x11C8
		x"FD",x"87",x"E4",x"20",x"00",x"01",x"14",x"01", -- 0x11D0
		x"15",x"FE",x"20",x"00",x"01",x"14",x"01",x"15", -- 0x11D8
		x"FE",x"FD",x"87",x"E4",x"20",x"00",x"01",x"14", -- 0x11E0
		x"01",x"15",x"10",x"22",x"FE",x"20",x"00",x"01", -- 0x11E8
		x"14",x"01",x"15",x"FE",x"FD",x"87",x"E5",x"20", -- 0x11F0
		x"00",x"01",x"14",x"01",x"15",x"28",x"00",x"FE", -- 0x11F8
		x"20",x"00",x"01",x"14",x"01",x"15",x"FE",x"FD", -- 0x1200
		x"87",x"E5",x"20",x"01",x"20",x"02",x"01",x"14", -- 0x1208
		x"01",x"15",x"04",x"01",x"FE",x"01",x"14",x"01", -- 0x1210
		x"15",x"20",x"01",x"20",x"02",x"04",x"40",x"FE", -- 0x1218
		x"FD",x"87",x"E5",x"01",x"14",x"01",x"15",x"20", -- 0x1220
		x"01",x"20",x"02",x"23",x"EA",x"04",x"01",x"FE", -- 0x1228
		x"20",x"01",x"20",x"02",x"01",x"14",x"01",x"15", -- 0x1230
		x"04",x"40",x"FE",x"FD",x"88",x"E5",x"00",x"12", -- 0x1238
		x"00",x"13",x"20",x"01",x"20",x"02",x"04",x"02", -- 0x1240
		x"FE",x"00",x"12",x"00",x"13",x"20",x"01",x"20", -- 0x1248
		x"02",x"04",x"40",x"FE",x"FD",x"88",x"E5",x"00", -- 0x1250
		x"12",x"00",x"13",x"20",x"01",x"20",x"02",x"10", -- 0x1258
		x"22",x"04",x"02",x"FE",x"00",x"12",x"00",x"13", -- 0x1260
		x"20",x"01",x"20",x"02",x"23",x"F3",x"04",x"40", -- 0x1268
		x"FE",x"FD",x"88",x"E5",x"00",x"12",x"00",x"13", -- 0x1270
		x"20",x"1A",x"20",x"1B",x"04",x"02",x"FE",x"00", -- 0x1278
		x"12",x"00",x"13",x"20",x"1A",x"20",x"1B",x"04", -- 0x1280
		x"40",x"FE",x"FD",x"86",x"E5",x"00",x"12",x"00", -- 0x1288
		x"13",x"20",x"1A",x"20",x"1B",x"28",x"00",x"04", -- 0x1290
		x"02",x"FE",x"00",x"12",x"00",x"13",x"20",x"1A", -- 0x1298
		x"20",x"1B",x"04",x"40",x"FE",x"FD",x"87",x"E5", -- 0x12A0
		x"00",x"12",x"00",x"13",x"20",x"1A",x"20",x"1B", -- 0x12A8
		x"04",x"02",x"FE",x"00",x"12",x"00",x"13",x"20", -- 0x12B0
		x"1A",x"20",x"1B",x"04",x"40",x"FE",x"FD",x"86", -- 0x12B8
		x"E4",x"00",x"12",x"00",x"13",x"20",x"1A",x"20", -- 0x12C0
		x"1B",x"FE",x"FE",x"FD",x"09",x"00",x"FD",x"FC", -- 0x12C8
		x"FF",x"80",x"C0",x"FE",x"FE",x"FD",x"86",x"C0", -- 0x12D0
		x"20",x"1A",x"20",x"1B",x"FE",x"20",x"1A",x"20", -- 0x12D8
		x"1B",x"FE",x"FD",x"86",x"C0",x"20",x"1A",x"20", -- 0x12E0
		x"1B",x"28",x"00",x"FE",x"20",x"1A",x"20",x"1B", -- 0x12E8
		x"FE",x"FD",x"86",x"C0",x"20",x"1A",x"20",x"1B", -- 0x12F0
		x"FE",x"20",x"1A",x"20",x"1B",x"10",x"65",x"FE", -- 0x12F8
		x"FD",x"86",x"C0",x"20",x"1A",x"20",x"1B",x"FE", -- 0x1300
		x"20",x"1A",x"20",x"1B",x"FE",x"FD",x"86",x"C0", -- 0x1308
		x"23",x"CC",x"FE",x"20",x"00",x"FE",x"FD",x"86", -- 0x1310
		x"C0",x"20",x"00",x"FE",x"20",x"00",x"10",x"63", -- 0x1318
		x"FE",x"FD",x"86",x"C0",x"20",x"00",x"FE",x"20", -- 0x1320
		x"00",x"10",x"66",x"FE",x"FD",x"87",x"C0",x"20", -- 0x1328
		x"00",x"FE",x"20",x"00",x"FE",x"FD",x"87",x"C0", -- 0x1330
		x"20",x"00",x"FE",x"10",x"64",x"FE",x"FD",x"87", -- 0x1338
		x"C0",x"20",x"01",x"20",x"02",x"FE",x"20",x"01", -- 0x1340
		x"20",x"02",x"FE",x"FD",x"86",x"C0",x"20",x"01", -- 0x1348
		x"20",x"02",x"28",x"00",x"FE",x"20",x"01",x"20", -- 0x1350
		x"02",x"FE",x"FD",x"86",x"C0",x"20",x"01",x"20", -- 0x1358
		x"02",x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x1360
		x"84",x"C0",x"20",x"01",x"20",x"02",x"FE",x"FE", -- 0x1368
		x"FD",x"FC",x"FF",x"80",x"C0",x"FE",x"FE",x"FD", -- 0x1370
		x"85",x"E4",x"00",x"16",x"00",x"17",x"FE",x"00", -- 0x1378
		x"16",x"00",x"17",x"10",x"24",x"FE",x"FD",x"85", -- 0x1380
		x"E4",x"00",x"16",x"00",x"17",x"23",x"C5",x"FE", -- 0x1388
		x"00",x"16",x"00",x"17",x"FE",x"FD",x"85",x"E4", -- 0x1390
		x"00",x"16",x"00",x"17",x"20",x"00",x"FE",x"00", -- 0x1398
		x"16",x"00",x"17",x"20",x"00",x"FE",x"FD",x"85", -- 0x13A0
		x"E4",x"00",x"16",x"00",x"17",x"20",x"00",x"10", -- 0x13A8
		x"21",x"FE",x"00",x"16",x"00",x"17",x"20",x"00", -- 0x13B0
		x"FE",x"FD",x"85",x"E5",x"00",x"18",x"00",x"19", -- 0x13B8
		x"20",x"00",x"28",x"00",x"FE",x"00",x"18",x"00", -- 0x13C0
		x"19",x"20",x"00",x"FE",x"FD",x"85",x"E5",x"00", -- 0x13C8
		x"18",x"00",x"19",x"20",x"00",x"FE",x"00",x"18", -- 0x13D0
		x"00",x"19",x"20",x"1E",x"20",x"1F",x"FE",x"FD", -- 0x13D8
		x"86",x"E5",x"00",x"18",x"00",x"19",x"20",x"1E", -- 0x13E0
		x"20",x"1F",x"23",x"CE",x"FE",x"00",x"18",x"00", -- 0x13E8
		x"19",x"20",x"1E",x"20",x"1F",x"FE",x"FD",x"86", -- 0x13F0
		x"E5",x"04",x"03",x"20",x"1E",x"20",x"1F",x"FE", -- 0x13F8
		x"20",x"1E",x"20",x"1F",x"FE",x"04",x"40",x"FD", -- 0x1400
		x"86",x"E5",x"04",x"03",x"20",x"1E",x"20",x"1F", -- 0x1408
		x"10",x"21",x"FE",x"23",x"D7",x"20",x"1E",x"20", -- 0x1410
		x"1F",x"FE",x"04",x"40",x"FD",x"86",x"E5",x"04", -- 0x1418
		x"03",x"20",x"01",x"20",x"02",x"FE",x"20",x"01", -- 0x1420
		x"20",x"02",x"FE",x"04",x"40",x"FD",x"85",x"E5", -- 0x1428
		x"04",x"03",x"20",x"01",x"20",x"02",x"28",x"00", -- 0x1430
		x"FE",x"20",x"01",x"20",x"02",x"FE",x"04",x"40", -- 0x1438
		x"FD",x"85",x"E5",x"04",x"03",x"20",x"01",x"20", -- 0x1440
		x"02",x"FE",x"20",x"01",x"20",x"02",x"FE",x"04", -- 0x1448
		x"40",x"FD",x"84",x"E2",x"04",x"03",x"20",x"01", -- 0x1450
		x"20",x"02",x"FE",x"FE",x"04",x"40",x"FD",x"FC", -- 0x1458
		x"FF",x"80",x"C0",x"FE",x"FE",x"FD",x"85",x"D4", -- 0x1460
		x"00",x"10",x"00",x"11",x"20",x"00",x"FE",x"00", -- 0x1468
		x"10",x"00",x"11",x"20",x"00",x"FE",x"FD",x"85", -- 0x1470
		x"D4",x"00",x"10",x"00",x"11",x"20",x"00",x"23", -- 0x1478
		x"D0",x"FE",x"00",x"10",x"00",x"11",x"20",x"00", -- 0x1480
		x"FE",x"FD",x"85",x"D4",x"00",x"10",x"00",x"11", -- 0x1488
		x"20",x"00",x"FE",x"00",x"10",x"00",x"11",x"20", -- 0x1490
		x"1A",x"20",x"1B",x"FE",x"FD",x"85",x"D4",x"00", -- 0x1498
		x"12",x"00",x"13",x"20",x"1A",x"20",x"1B",x"10", -- 0x14A0
		x"20",x"FE",x"00",x"12",x"00",x"13",x"20",x"1A", -- 0x14A8
		x"20",x"1B",x"FE",x"FD",x"85",x"D5",x"00",x"12", -- 0x14B0
		x"00",x"13",x"20",x"1A",x"20",x"1B",x"28",x"00", -- 0x14B8
		x"FE",x"00",x"12",x"00",x"13",x"20",x"1A",x"20", -- 0x14C0
		x"1B",x"FE",x"FD",x"85",x"D5",x"00",x"12",x"00", -- 0x14C8
		x"13",x"20",x"1A",x"20",x"1B",x"FE",x"00",x"12", -- 0x14D0
		x"00",x"13",x"20",x"1A",x"20",x"1B",x"FE",x"FD", -- 0x14D8
		x"86",x"D5",x"20",x"18",x"20",x"19",x"00",x"03", -- 0x14E0
		x"00",x"04",x"03",x"E1",x"FE",x"20",x"18",x"20", -- 0x14E8
		x"19",x"00",x"03",x"00",x"04",x"FE",x"FD",x"86", -- 0x14F0
		x"D5",x"20",x"18",x"20",x"19",x"00",x"03",x"00", -- 0x14F8
		x"04",x"FE",x"20",x"18",x"20",x"19",x"00",x"03", -- 0x1500
		x"00",x"04",x"FE",x"FD",x"86",x"D5",x"20",x"18", -- 0x1508
		x"20",x"19",x"00",x"03",x"00",x"04",x"10",x"20", -- 0x1510
		x"FE",x"20",x"18",x"20",x"19",x"00",x"03",x"00", -- 0x1518
		x"04",x"03",x"EA",x"FE",x"FD",x"87",x"D5",x"20", -- 0x1520
		x"1E",x"20",x"1F",x"00",x"14",x"00",x"15",x"FE", -- 0x1528
		x"20",x"1E",x"20",x"1F",x"00",x"14",x"00",x"15", -- 0x1530
		x"FE",x"FD",x"86",x"D5",x"20",x"1E",x"20",x"1F", -- 0x1538
		x"00",x"14",x"00",x"15",x"28",x"00",x"FE",x"20", -- 0x1540
		x"1E",x"20",x"1F",x"00",x"14",x"00",x"15",x"FE", -- 0x1548
		x"FD",x"86",x"D5",x"20",x"1E",x"20",x"1F",x"00", -- 0x1550
		x"14",x"00",x"15",x"FE",x"20",x"1E",x"20",x"1F", -- 0x1558
		x"00",x"14",x"00",x"15",x"FE",x"FD",x"85",x"D4", -- 0x1560
		x"20",x"1E",x"20",x"1F",x"00",x"14",x"00",x"15", -- 0x1568
		x"FE",x"FE",x"FD",x"FC",x"FF",x"80",x"C0",x"FE", -- 0x1570
		x"FE",x"FD",x"87",x"E5",x"01",x"03",x"01",x"04", -- 0x1578
		x"20",x"00",x"FE",x"01",x"03",x"01",x"04",x"20", -- 0x1580
		x"00",x"FE",x"FD",x"87",x"E5",x"01",x"03",x"01", -- 0x1588
		x"04",x"20",x"00",x"23",x"E3",x"FE",x"01",x"03", -- 0x1590
		x"01",x"04",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x1598
		x"87",x"E6",x"01",x"03",x"01",x"04",x"20",x"01", -- 0x15A0
		x"20",x"02",x"FE",x"01",x"03",x"01",x"04",x"20", -- 0x15A8
		x"01",x"20",x"02",x"FE",x"FD",x"87",x"E6",x"01", -- 0x15B0
		x"12",x"01",x"13",x"20",x"01",x"20",x"02",x"10", -- 0x15B8
		x"22",x"FE",x"01",x"12",x"01",x"13",x"20",x"01", -- 0x15C0
		x"20",x"02",x"FE",x"FD",x"87",x"E6",x"01",x"12", -- 0x15C8
		x"01",x"13",x"20",x"01",x"20",x"02",x"28",x"00", -- 0x15D0
		x"FE",x"01",x"12",x"01",x"13",x"20",x"01",x"20", -- 0x15D8
		x"02",x"FE",x"FD",x"88",x"E6",x"01",x"12",x"01", -- 0x15E0
		x"13",x"20",x"01",x"20",x"02",x"FE",x"01",x"12", -- 0x15E8
		x"01",x"13",x"20",x"1C",x"20",x"1D",x"FE",x"FD", -- 0x15F0
		x"88",x"E6",x"01",x"12",x"01",x"13",x"20",x"1C", -- 0x15F8
		x"20",x"1D",x"23",x"EC",x"FE",x"01",x"12",x"01", -- 0x1600
		x"13",x"20",x"1C",x"20",x"1D",x"FE",x"FD",x"88", -- 0x1608
		x"E6",x"00",x"16",x"00",x"17",x"20",x"1C",x"20", -- 0x1610
		x"1D",x"FE",x"00",x"16",x"00",x"17",x"20",x"1C", -- 0x1618
		x"20",x"1D",x"FE",x"FD",x"88",x"E6",x"00",x"16", -- 0x1620
		x"00",x"17",x"20",x"1C",x"20",x"1D",x"10",x"22", -- 0x1628
		x"FE",x"00",x"16",x"00",x"17",x"20",x"1C",x"20", -- 0x1630
		x"1D",x"23",x"F5",x"FE",x"FD",x"88",x"E7",x"00", -- 0x1638
		x"16",x"00",x"17",x"20",x"1C",x"20",x"1D",x"FE", -- 0x1640
		x"00",x"16",x"00",x"17",x"20",x"1C",x"20",x"1D", -- 0x1648
		x"FE",x"FD",x"88",x"E7",x"00",x"16",x"00",x"17", -- 0x1650
		x"20",x"1E",x"20",x"1F",x"28",x"00",x"FE",x"00", -- 0x1658
		x"16",x"00",x"17",x"20",x"1E",x"20",x"1F",x"FE", -- 0x1660
		x"FD",x"87",x"E6",x"00",x"16",x"00",x"17",x"20", -- 0x1668
		x"1E",x"20",x"1F",x"FE",x"00",x"16",x"00",x"17", -- 0x1670
		x"20",x"1E",x"20",x"1F",x"FE",x"FD",x"85",x"E3", -- 0x1678
		x"00",x"16",x"00",x"17",x"20",x"1E",x"20",x"1F", -- 0x1680
		x"FE",x"FE",x"FD",x"FC",x"FF",x"80",x"C0",x"FE", -- 0x1688
		x"FE",x"FD",x"85",x"C0",x"23",x"E6",x"FE",x"20", -- 0x1690
		x"01",x"20",x"02",x"FE",x"FD",x"85",x"C0",x"20", -- 0x1698
		x"01",x"20",x"02",x"FE",x"20",x"01",x"20",x"02", -- 0x16A0
		x"10",x"65",x"FE",x"FD",x"85",x"C0",x"20",x"01", -- 0x16A8
		x"20",x"02",x"FE",x"20",x"01",x"20",x"02",x"FE", -- 0x16B0
		x"FD",x"86",x"C0",x"20",x"01",x"20",x"02",x"10", -- 0x16B8
		x"64",x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD", -- 0x16C0
		x"86",x"C0",x"20",x"01",x"20",x"02",x"FE",x"23", -- 0x16C8
		x"EF",x"FE",x"FD",x"86",x"C0",x"20",x"1A",x"20", -- 0x16D0
		x"1B",x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD", -- 0x16D8
		x"86",x"C0",x"20",x"1A",x"20",x"1B",x"10",x"62", -- 0x16E0
		x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD",x"85", -- 0x16E8
		x"C0",x"20",x"1A",x"20",x"1B",x"10",x"66",x"FE", -- 0x16F0
		x"20",x"1A",x"20",x"1B",x"FE",x"FD",x"85",x"C0", -- 0x16F8
		x"20",x"1A",x"20",x"1B",x"FE",x"10",x"63",x"FE", -- 0x1700
		x"FD",x"85",x"C0",x"20",x"00",x"FE",x"20",x"00", -- 0x1708
		x"FE",x"FD",x"84",x"C0",x"20",x"00",x"28",x"00", -- 0x1710
		x"FE",x"20",x"00",x"FE",x"FD",x"85",x"C0",x"20", -- 0x1718
		x"00",x"FE",x"20",x"00",x"FE",x"FD",x"84",x"C0", -- 0x1720
		x"20",x"00",x"FE",x"FE",x"FD",x"FC",x"FF",x"80", -- 0x1728
		x"C0",x"FE",x"FE",x"FD",x"86",x"E4",x"20",x"00", -- 0x1730
		x"04",x"03",x"FE",x"20",x"00",x"10",x"24",x"FE", -- 0x1738
		x"04",x"40",x"FD",x"86",x"E4",x"20",x"00",x"04", -- 0x1740
		x"03",x"23",x"C0",x"FE",x"20",x"01",x"20",x"02", -- 0x1748
		x"FE",x"04",x"40",x"FD",x"86",x"E5",x"20",x"01", -- 0x1750
		x"20",x"02",x"04",x"03",x"FE",x"20",x"01",x"20", -- 0x1758
		x"02",x"FE",x"04",x"40",x"FD",x"86",x"E5",x"20", -- 0x1760
		x"01",x"20",x"02",x"04",x"03",x"10",x"21",x"FE", -- 0x1768
		x"20",x"01",x"20",x"02",x"FE",x"04",x"40",x"FD", -- 0x1770
		x"87",x"E5",x"20",x"01",x"20",x"02",x"04",x"04", -- 0x1778
		x"28",x"00",x"FE",x"20",x"01",x"20",x"02",x"FE", -- 0x1780
		x"04",x"40",x"FD",x"87",x"E6",x"04",x"04",x"20", -- 0x1788
		x"1A",x"20",x"1B",x"FE",x"20",x"1A",x"20",x"1B", -- 0x1790
		x"FE",x"04",x"40",x"FD",x"87",x"E6",x"01",x"03", -- 0x1798
		x"01",x"04",x"20",x"1A",x"20",x"1B",x"23",x"C9", -- 0x17A0
		x"FE",x"01",x"03",x"01",x"04",x"20",x"1A",x"20", -- 0x17A8
		x"1B",x"FE",x"FD",x"87",x"E6",x"01",x"03",x"01", -- 0x17B0
		x"04",x"20",x"1A",x"20",x"1B",x"FE",x"01",x"03", -- 0x17B8
		x"01",x"04",x"20",x"1A",x"20",x"1B",x"FE",x"FD", -- 0x17C0
		x"88",x"E6",x"01",x"03",x"01",x"04",x"20",x"1A", -- 0x17C8
		x"20",x"1B",x"10",x"21",x"FE",x"01",x"03",x"01", -- 0x17D0
		x"04",x"20",x"1A",x"20",x"1B",x"23",x"D2",x"FE", -- 0x17D8
		x"FD",x"89",x"E6",x"01",x"12",x"01",x"13",x"20", -- 0x17E0
		x"1E",x"20",x"1F",x"FE",x"01",x"12",x"01",x"13", -- 0x17E8
		x"20",x"1E",x"20",x"1F",x"FE",x"FD",x"87",x"E6", -- 0x17F0
		x"01",x"12",x"01",x"13",x"20",x"1E",x"20",x"1F", -- 0x17F8
		x"28",x"00",x"FE",x"01",x"12",x"01",x"13",x"20", -- 0x1800
		x"1E",x"20",x"1F",x"FE",x"FD",x"88",x"E5",x"01", -- 0x1808
		x"12",x"01",x"13",x"20",x"1E",x"20",x"1F",x"FE", -- 0x1810
		x"01",x"12",x"01",x"13",x"20",x"1E",x"20",x"1F", -- 0x1818
		x"FE",x"FD",x"86",x"E3",x"01",x"12",x"01",x"13", -- 0x1820
		x"20",x"1E",x"20",x"1F",x"FE",x"FE",x"FD",x"FC", -- 0x1828
		x"FF",x"80",x"C0",x"FE",x"FE",x"FD",x"89",x"E5", -- 0x1830
		x"01",x"03",x"01",x"04",x"20",x"12",x"20",x"13", -- 0x1838
		x"FE",x"01",x"03",x"01",x"04",x"20",x"12",x"20", -- 0x1840
		x"13",x"FE",x"FD",x"89",x"E5",x"23",x"D3",x"01", -- 0x1848
		x"03",x"01",x"04",x"20",x"12",x"20",x"13",x"FE", -- 0x1850
		x"01",x"03",x"01",x"04",x"20",x"12",x"20",x"13", -- 0x1858
		x"FE",x"FD",x"89",x"E5",x"01",x"03",x"01",x"04", -- 0x1860
		x"20",x"12",x"20",x"13",x"FE",x"01",x"03",x"01", -- 0x1868
		x"04",x"20",x"12",x"20",x"13",x"FE",x"FD",x"89", -- 0x1870
		x"E6",x"01",x"12",x"01",x"13",x"20",x"10",x"20", -- 0x1878
		x"11",x"10",x"20",x"FE",x"01",x"12",x"01",x"13", -- 0x1880
		x"20",x"10",x"20",x"11",x"FE",x"FD",x"89",x"E6", -- 0x1888
		x"28",x"00",x"01",x"12",x"01",x"13",x"20",x"10", -- 0x1890
		x"20",x"11",x"FE",x"01",x"12",x"01",x"13",x"20", -- 0x1898
		x"10",x"20",x"11",x"FE",x"FD",x"89",x"C6",x"01", -- 0x18A0
		x"12",x"01",x"13",x"20",x"10",x"20",x"11",x"FE", -- 0x18A8
		x"01",x"12",x"01",x"13",x"20",x"10",x"20",x"11", -- 0x18B0
		x"FE",x"FD",x"8A",x"C6",x"20",x"1C",x"20",x"1D", -- 0x18B8
		x"04",x"03",x"23",x"E4",x"FE",x"20",x"1C",x"20", -- 0x18C0
		x"1D",x"FE",x"04",x"40",x"FD",x"8A",x"C6",x"20", -- 0x18C8
		x"1C",x"20",x"1D",x"04",x"03",x"FE",x"20",x"1C", -- 0x18D0
		x"20",x"1D",x"FE",x"04",x"40",x"FD",x"8A",x"C6", -- 0x18D8
		x"20",x"1E",x"20",x"1F",x"04",x"03",x"10",x"20", -- 0x18E0
		x"FE",x"20",x"1E",x"20",x"1F",x"23",x"ED",x"FE", -- 0x18E8
		x"04",x"40",x"FD",x"8A",x"C6",x"20",x"1E",x"20", -- 0x18F0
		x"1F",x"04",x"03",x"FE",x"20",x"1E",x"20",x"1F", -- 0x18F8
		x"FE",x"04",x"40",x"FD",x"89",x"C6",x"20",x"1E", -- 0x1900
		x"20",x"1F",x"04",x"03",x"28",x"00",x"FE",x"20", -- 0x1908
		x"1E",x"20",x"1F",x"FE",x"04",x"40",x"FD",x"8A", -- 0x1910
		x"C6",x"20",x"1E",x"20",x"1F",x"04",x"03",x"FE", -- 0x1918
		x"20",x"1E",x"20",x"1F",x"FE",x"04",x"40",x"FD", -- 0x1920
		x"89",x"C6",x"20",x"1E",x"20",x"1F",x"04",x"03", -- 0x1928
		x"FE",x"FE",x"04",x"40",x"FD",x"FC",x"FF",x"80", -- 0x1930
		x"C0",x"FE",x"FE",x"FD",x"89",x"C6",x"20",x"00", -- 0x1938
		x"04",x"04",x"01",x"03",x"01",x"04",x"FE",x"01", -- 0x1940
		x"03",x"01",x"04",x"20",x"00",x"FE",x"04",x"40", -- 0x1948
		x"FD",x"89",x"C6",x"20",x"00",x"04",x"04",x"01", -- 0x1950
		x"03",x"01",x"04",x"23",x"EE",x"FE",x"01",x"03", -- 0x1958
		x"01",x"04",x"20",x"00",x"FE",x"04",x"40",x"FD", -- 0x1960
		x"89",x"C6",x"20",x"01",x"20",x"02",x"04",x"04", -- 0x1968
		x"01",x"03",x"01",x"04",x"FE",x"01",x"03",x"01", -- 0x1970
		x"04",x"20",x"01",x"20",x"02",x"FE",x"04",x"40", -- 0x1978
		x"FD",x"8A",x"C6",x"20",x"1A",x"20",x"1B",x"04", -- 0x1980
		x"04",x"01",x"03",x"01",x"04",x"10",x"22",x"FE", -- 0x1988
		x"01",x"03",x"01",x"04",x"20",x"1A",x"20",x"1B", -- 0x1990
		x"FE",x"04",x"40",x"FD",x"8A",x"C6",x"04",x"04", -- 0x1998
		x"28",x"00",x"20",x"1A",x"20",x"1B",x"00",x"12", -- 0x19A0
		x"00",x"13",x"FE",x"20",x"1A",x"20",x"1B",x"00", -- 0x19A8
		x"12",x"00",x"13",x"FE",x"04",x"40",x"FD",x"8A", -- 0x19B0
		x"C7",x"04",x"04",x"20",x"1A",x"20",x"1B",x"00", -- 0x19B8
		x"12",x"00",x"13",x"FE",x"00",x"12",x"00",x"13", -- 0x19C0
		x"20",x"1A",x"20",x"1B",x"FE",x"04",x"40",x"FD", -- 0x19C8
		x"8A",x"E7",x"20",x"1C",x"20",x"1D",x"04",x"05", -- 0x19D0
		x"00",x"12",x"00",x"13",x"23",x"F7",x"FE",x"00", -- 0x19D8
		x"12",x"00",x"13",x"20",x"1C",x"20",x"1D",x"FE", -- 0x19E0
		x"04",x"40",x"FD",x"8A",x"E7",x"04",x"05",x"00", -- 0x19E8
		x"14",x"00",x"15",x"20",x"1C",x"20",x"1D",x"FE", -- 0x19F0
		x"00",x"14",x"00",x"15",x"20",x"1C",x"20",x"1D", -- 0x19F8
		x"FE",x"04",x"40",x"FD",x"8B",x"E7",x"00",x"18", -- 0x1A00
		x"00",x"19",x"20",x"1C",x"20",x"1D",x"10",x"22", -- 0x1A08
		x"FE",x"00",x"18",x"00",x"19",x"20",x"1C",x"20", -- 0x1A10
		x"1D",x"FE",x"23",x"D0",x"FD",x"8B",x"E7",x"20", -- 0x1A18
		x"1E",x"20",x"1F",x"00",x"18",x"00",x"19",x"FE", -- 0x1A20
		x"20",x"1E",x"20",x"1F",x"00",x"16",x"00",x"17", -- 0x1A28
		x"FE",x"FD",x"89",x"E8",x"20",x"1E",x"20",x"1F", -- 0x1A30
		x"28",x"00",x"00",x"16",x"00",x"17",x"FE",x"20", -- 0x1A38
		x"1E",x"20",x"1F",x"00",x"16",x"00",x"17",x"FE", -- 0x1A40
		x"FD",x"8A",x"E8",x"20",x"1E",x"20",x"1F",x"00", -- 0x1A48
		x"16",x"00",x"17",x"FE",x"20",x"1E",x"20",x"1F", -- 0x1A50
		x"00",x"16",x"00",x"17",x"FE",x"FD",x"8A",x"E8", -- 0x1A58
		x"20",x"1E",x"20",x"1F",x"00",x"16",x"00",x"17", -- 0x1A60
		x"FE",x"FE",x"FD",x"29",x"01",x"FD",x"FC",x"FF", -- 0x1A68
		x"80",x"C0",x"FE",x"FE",x"FD",x"84",x"C0",x"10", -- 0x1A70
		x"60",x"FE",x"20",x"00",x"FE",x"FD",x"84",x"C0", -- 0x1A78
		x"20",x"00",x"10",x"61",x"FE",x"20",x"00",x"FE", -- 0x1A80
		x"FD",x"84",x"C0",x"20",x"00",x"FE",x"23",x"E1", -- 0x1A88
		x"FE",x"FD",x"84",x"C0",x"20",x"01",x"20",x"02", -- 0x1A90
		x"FE",x"20",x"01",x"20",x"02",x"FE",x"FD",x"83", -- 0x1A98
		x"C0",x"20",x"01",x"20",x"02",x"FE",x"20",x"01", -- 0x1AA0
		x"20",x"02",x"23",x"CA",x"FE",x"FD",x"83",x"C0", -- 0x1AA8
		x"20",x"01",x"20",x"02",x"FE",x"20",x"01",x"20", -- 0x1AB0
		x"02",x"23",x"D3",x"FE",x"FD",x"84",x"C0",x"20", -- 0x1AB8
		x"01",x"20",x"02",x"FE",x"20",x"01",x"20",x"02", -- 0x1AC0
		x"FE",x"FD",x"85",x"C0",x"20",x"01",x"20",x"02", -- 0x1AC8
		x"FE",x"10",x"63",x"FE",x"FD",x"85",x"C0",x"20", -- 0x1AD0
		x"1A",x"20",x"1B",x"FE",x"20",x"1A",x"20",x"1B", -- 0x1AD8
		x"FE",x"FD",x"84",x"C0",x"20",x"1A",x"20",x"1B", -- 0x1AE0
		x"10",x"20",x"FE",x"20",x"1A",x"20",x"1B",x"FE", -- 0x1AE8
		x"FD",x"83",x"C0",x"20",x"1A",x"20",x"1B",x"28", -- 0x1AF0
		x"00",x"FE",x"20",x"1A",x"20",x"1B",x"FE",x"FD", -- 0x1AF8
		x"84",x"C0",x"20",x"1A",x"20",x"1B",x"FE",x"20", -- 0x1B00
		x"1A",x"20",x"1B",x"FE",x"FD",x"83",x"C0",x"20", -- 0x1B08
		x"1A",x"20",x"1B",x"FE",x"FE",x"FD",x"FC",x"FF", -- 0x1B10
		x"0E",x"51",x"50",x"AF",x"C1",x"D0",x"73",x"52", -- 0x1B18
		x"98",x"05",x"26",x"84",x"80",x"26",x"05",x"A0", -- 0x1B20
		x"14",x"44",x"88",x"D7",x"00",x"35",x"00",x"80", -- 0x1B28
		x"00",x"01",x"9C",x"40",x"04",x"2F",x"37",x"48", -- 0x1B30
		x"34",x"DD",x"22",x"99",x"C5",x"B7",x"00",x"04", -- 0x1B38
		x"24",x"21",x"02",x"6A",x"85",x"3F",x"41",x"2E", -- 0x1B40
		x"50",x"E0",x"80",x"61",x"C0",x"4B",x"79",x"1C", -- 0x1B48
		x"58",x"F7",x"86",x"1B",x"E8",x"00",x"07",x"8B", -- 0x1B50
		x"72",x"67",x"09",x"03",x"A8",x"75",x"C0",x"EC", -- 0x1B58
		x"C0",x"EC",x"05",x"66",x"A8",x"D6",x"18",x"6D", -- 0x1B60
		x"C4",x"1C",x"54",x"9E",x"A0",x"28",x"08",x"92", -- 0x1B68
		x"98",x"38",x"A5",x"C5",x"40",x"EA",x"C8",x"43", -- 0x1B70
		x"12",x"01",x"61",x"0A",x"50",x"04",x"2A",x"0C", -- 0x1B78
		x"06",x"CA",x"69",x"1C",x"04",x"46",x"01",x"9F", -- 0x1B80
		x"01",x"63",x"80",x"20",x"00",x"C2",x"10",x"51", -- 0x1B88
		x"40",x"03",x"42",x"35",x"00",x"25",x"49",x"0E", -- 0x1B90
		x"FC",x"00",x"79",x"E0",x"04",x"30",x"A4",x"52", -- 0x1B98
		x"20",x"41",x"80",x"4D",x"C5",x"31",x"01",x"8C", -- 0x1BA0
		x"1B",x"E4",x"01",x"07",x"80",x"4A",x"41",x"A8", -- 0x1BA8
		x"14",x"A3",x"20",x"D4",x"A0",x"02",x"C2",x"5C", -- 0x1BB0
		x"16",x"91",x"30",x"25",x"40",x"02",x"19",x"CE", -- 0x1BB8
		x"30",x"26",x"C2",x"A7",x"8A",x"CC",x"19",x"14", -- 0x1BC0
		x"61",x"C5",x"3D",x"C5",x"0C",x"B5",x"43",x"03", -- 0x1BC8
		x"12",x"0E",x"11",x"E2",x"90",x"98",x"06",x"A1", -- 0x1BD0
		x"94",x"6C",x"41",x"2E",x"EA",x"24",x"28",x"98", -- 0x1BD8
		x"04",x"AF",x"40",x"2E",x"04",x"56",x"01",x"4A", -- 0x1BE0
		x"D4",x"69",x"28",x"5D",x"C4",x"C3",x"AD",x"06", -- 0x1BE8
		x"00",x"AA",x"44",x"29",x"4E",x"78",x"80",x"9E", -- 0x1BF0
		x"91",x"08",x"44",x"52",x"48",x"42",x"44",x"71", -- 0x1BF8
		x"40",x"04",x"A0",x"65",x"2C",x"F0",x"C1",x"01", -- 0x1C00
		x"02",x"64",x"78",x"06",x"49",x"24",x"23",x"40", -- 0x1C08
		x"C8",x"26",x"0B",x"82",x"29",x"05",x"A3",x"EB", -- 0x1C10
		x"45",x"05",x"95",x"72",x"4E",x"27",x"64",x"00", -- 0x1C18
		x"00",x"DC",x"04",x"44",x"A4",x"B5",x"16",x"01", -- 0x1C20
		x"45",x"40",x"A4",x"06",x"08",x"24",x"0A",x"20", -- 0x1C28
		x"4D",x"C4",x"88",x"07",x"08",x"A3",x"52",x"08", -- 0x1C30
		x"21",x"FC",x"03",x"09",x"9C",x"2D",x"40",x"08", -- 0x1C38
		x"03",x"A8",x"00",x"49",x"0F",x"32",x"0B",x"22", -- 0x1C40
		x"39",x"B0",x"98",x"88",x"79",x"13",x"22",x"00", -- 0x1C48
		x"1C",x"E8",x"44",x"60",x"81",x"DD",x"10",x"89", -- 0x1C50
		x"1C",x"96",x"1F",x"02",x"C1",x"6B",x"14",x"10", -- 0x1C58
		x"58",x"61",x"05",x"83",x"08",x"42",x"62",x"18", -- 0x1C60
		x"1A",x"40",x"01",x"23",x"3A",x"03",x"C4",x"03", -- 0x1C68
		x"44",x"0F",x"14",x"74",x"38",x"ED",x"00",x"AC", -- 0x1C70
		x"3C",x"01",x"65",x"CB",x"09",x"89",x"07",x"3A", -- 0x1C78
		x"E8",x"60",x"50",x"16",x"8A",x"58",x"10",x"23", -- 0x1C80
		x"1C",x"50",x"92",x"46",x"60",x"64",x"2C",x"3C", -- 0x1C88
		x"20",x"11",x"A6",x"34",x"A2",x"11",x"00",x"99", -- 0x1C90
		x"30",x"E0",x"09",x"C3",x"01",x"AB",x"C0",x"42", -- 0x1C98
		x"01",x"82",x"22",x"AB",x"49",x"04",x"48",x"47", -- 0x1CA0
		x"82",x"3B",x"A0",x"02",x"A0",x"1F",x"91",x"76", -- 0x1CA8
		x"70",x"B1",x"22",x"48",x"00",x"C4",x"4A",x"12", -- 0x1CB0
		x"0E",x"23",x"05",x"B9",x"18",x"CF",x"65",x"C3", -- 0x1CB8
		x"01",x"04",x"61",x"EE",x"5A",x"BC",x"08",x"05", -- 0x1CC0
		x"B8",x"34",x"F9",x"70",x"D1",x"63",x"6E",x"B1", -- 0x1CC8
		x"00",x"41",x"46",x"C2",x"40",x"37",x"44",x"CA", -- 0x1CD0
		x"08",x"26",x"9F",x"AB",x"01",x"10",x"CC",x"02", -- 0x1CD8
		x"10",x"E6",x"01",x"5A",x"21",x"CB",x"33",x"09", -- 0x1CE0
		x"0F",x"D2",x"9C",x"0E",x"C2",x"53",x"7D",x"00", -- 0x1CE8
		x"10",x"C8",x"92",x"F1",x"11",x"B1",x"49",x"82", -- 0x1CF0
		x"00",x"F4",x"40",x"5C",x"28",x"32",x"61",x"02", -- 0x1CF8
		x"40",x"F0",x"91",x"86",x"69",x"31",x"EA",x"80", -- 0x1D00
		x"B0",x"8A",x"18",x"C2",x"C6",x"A4",x"10",x"06", -- 0x1D08
		x"00",x"B4",x"C4",x"C0",x"51",x"D2",x"84",x"23", -- 0x1D10
		x"0C",x"8C",x"93",x"04",x"01",x"05",x"A8",x"51", -- 0x1D18
		x"60",x"73",x"96",x"8F",x"40",x"1F",x"00",x"9D", -- 0x1D20
		x"99",x"6B",x"96",x"A8",x"80",x"4A",x"68",x"08", -- 0x1D28
		x"12",x"0B",x"31",x"D0",x"00",x"6A",x"14",x"1A", -- 0x1D30
		x"23",x"15",x"09",x"A6",x"58",x"2C",x"25",x"59", -- 0x1D38
		x"50",x"93",x"44",x"00",x"00",x"22",x"06",x"C3", -- 0x1D40
		x"DA",x"D0",x"29",x"A8",x"7A",x"03",x"BC",x"44", -- 0x1D48
		x"21",x"08",x"4A",x"09",x"C0",x"C0",x"AB",x"63", -- 0x1D50
		x"44",x"5C",x"26",x"72",x"ED",x"EC",x"20",x"10", -- 0x1D58
		x"00",x"59",x"50",x"9C",x"76",x"F7",x"B0",x"A3", -- 0x1D60
		x"80",x"18",x"08",x"81",x"15",x"10",x"FA",x"07", -- 0x1D68
		x"C0",x"41",x"0B",x"D6",x"4C",x"86",x"14",x"23", -- 0x1D70
		x"CE",x"04",x"36",x"70",x"01",x"88",x"00",x"10", -- 0x1D78
		x"74",x"43",x"1C",x"61",x"25",x"01",x"81",x"46", -- 0x1D80
		x"3F",x"28",x"FC",x"11",x"C8",x"4A",x"29",x"14", -- 0x1D88
		x"50",x"E4",x"FC",x"0A",x"14",x"40",x"80",x"88", -- 0x1D90
		x"71",x"09",x"0E",x"8A",x"56",x"21",x"3A",x"0A", -- 0x1D98
		x"08",x"56",x"14",x"F8",x"05",x"31",x"94",x"06", -- 0x1DA0
		x"B4",x"03",x"4B",x"4B",x"04",x"26",x"87",x"2D", -- 0x1DA8
		x"80",x"BB",x"11",x"C8",x"A6",x"A6",x"02",x"21", -- 0x1DB0
		x"A0",x"F9",x"83",x"A1",x"04",x"02",x"37",x"C8", -- 0x1DB8
		x"08",x"62",x"42",x"B0",x"83",x"A9",x"0A",x"31", -- 0x1DC0
		x"B6",x"C7",x"4A",x"A9",x"1A",x"93",x"58",x"15", -- 0x1DC8
		x"0E",x"66",x"2D",x"2C",x"34",x"35",x"91",x"B9", -- 0x1DD0
		x"85",x"20",x"12",x"84",x"4A",x"90",x"68",x"04", -- 0x1DD8
		x"18",x"10",x"A2",x"85",x"96",x"72",x"28",x"60", -- 0x1DE0
		x"A8",x"69",x"23",x"19",x"26",x"13",x"0F",x"B1", -- 0x1DE8
		x"40",x"25",x"11",x"90",x"01",x"52",x"13",x"C4", -- 0x1DF0
		x"D2",x"DE",x"00",x"89",x"60",x"69",x"88",x"21", -- 0x1DF8
		x"57",x"02",x"C3",x"2E",x"6E",x"81",x"64",x"5A", -- 0x1E00
		x"DE",x"9A",x"AC",x"93",x"24",x"C9",x"47",x"02", -- 0x1E08
		x"00",x"03",x"80",x"CD",x"18",x"8C",x"10",x"02", -- 0x1E10
		x"56",x"04",x"09",x"FD",x"88",x"42",x"17",x"04", -- 0x1E18
		x"04",x"BB",x"23",x"DA",x"3A",x"8A",x"03",x"99", -- 0x1E20
		x"3C",x"21",x"88",x"82",x"7A",x"0A",x"46",x"43", -- 0x1E28
		x"42",x"6C",x"82",x"02",x"4E",x"B6",x"82",x"60", -- 0x1E30
		x"6C",x"4C",x"24",x"CE",x"23",x"8E",x"01",x"91", -- 0x1E38
		x"C0",x"D8",x"D8",x"29",x"CB",x"90",x"66",x"20", -- 0x1E40
		x"AC",x"E0",x"E5",x"A3",x"DC",x"00",x"D2",x"02", -- 0x1E48
		x"0A",x"30",x"C1",x"40",x"B8",x"C4",x"40",x"E5", -- 0x1E50
		x"E4",x"C2",x"1D",x"21",x"A2",x"0A",x"23",x"91", -- 0x1E58
		x"14",x"A4",x"C4",x"00",x"10",x"AF",x"47",x"0A", -- 0x1E60
		x"93",x"72",x"02",x"A0",x"24",x"09",x"E0",x"0D", -- 0x1E68
		x"01",x"40",x"64",x"C9",x"10",x"08",x"32",x"A8", -- 0x1E70
		x"28",x"88",x"14",x"61",x"E1",x"E0",x"02",x"48", -- 0x1E78
		x"22",x"D6",x"87",x"A2",x"71",x"89",x"45",x"02", -- 0x1E80
		x"00",x"C8",x"91",x"21",x"1C",x"20",x"39",x"40", -- 0x1E88
		x"81",x"92",x"96",x"8D",x"09",x"71",x"17",x"6C", -- 0x1E90
		x"83",x"27",x"CC",x"94",x"A0",x"0A",x"2A",x"66", -- 0x1E98
		x"02",x"22",x"64",x"87",x"CA",x"12",x"B6",x"87", -- 0x1EA0
		x"30",x"81",x"41",x"E9",x"80",x"9A",x"54",x"57", -- 0x1EA8
		x"28",x"1D",x"A5",x"00",x"05",x"36",x"10",x"32", -- 0x1EB0
		x"28",x"A3",x"00",x"D0",x"CA",x"15",x"00",x"22", -- 0x1EB8
		x"02",x"98",x"30",x"8D",x"A6",x"C9",x"87",x"82", -- 0x1EC0
		x"83",x"8D",x"AA",x"4C",x"9C",x"A2",x"29",x"10", -- 0x1EC8
		x"50",x"05",x"18",x"80",x"D7",x"80",x"16",x"98", -- 0x1ED0
		x"9C",x"1C",x"1A",x"21",x"38",x"92",x"01",x"6F", -- 0x1ED8
		x"08",x"03",x"61",x"04",x"94",x"22",x"05",x"20", -- 0x1EE0
		x"06",x"F1",x"5F",x"B0",x"50",x"82",x"60",x"20", -- 0x1EE8
		x"0C",x"EB",x"48",x"07",x"A4",x"08",x"5E",x"04", -- 0x1EF0
		x"08",x"81",x"43",x"C8",x"28",x"81",x"4D",x"58", -- 0x1EF8
		x"25",x"E6",x"CC",x"60",x"7A",x"15",x"D3",x"A6", -- 0x1F00
		x"44",x"41",x"11",x"E6",x"2E",x"46",x"FB",x"C5", -- 0x1F08
		x"16",x"1D",x"5C",x"A2",x"0D",x"76",x"82",x"8A", -- 0x1F10
		x"2A",x"38",x"CD",x"5C",x"CE",x"89",x"A7",x"05", -- 0x1F18
		x"08",x"02",x"4F",x"88",x"88",x"3C",x"42",x"20", -- 0x1F20
		x"B0",x"18",x"42",x"C2",x"02",x"A3",x"CC",x"C2", -- 0x1F28
		x"10",x"10",x"09",x"D5",x"CE",x"84",x"28",x"1D", -- 0x1F30
		x"24",x"60",x"62",x"CE",x"14",x"4E",x"62",x"10", -- 0x1F38
		x"0E",x"0D",x"A5",x"00",x"32",x"68",x"60",x"00", -- 0x1F40
		x"80",x"70",x"00",x"18",x"BE",x"5B",x"68",x"61", -- 0x1F48
		x"46",x"31",x"D9",x"3D",x"06",x"09",x"61",x"39", -- 0x1F50
		x"50",x"07",x"C9",x"82",x"16",x"28",x"62",x"48", -- 0x1F58
		x"02",x"C8",x"A8",x"17",x"C2",x"61",x"28",x"98", -- 0x1F60
		x"00",x"81",x"9B",x"22",x"0C",x"44",x"38",x"22", -- 0x1F68
		x"48",x"E0",x"44",x"4D",x"05",x"10",x"26",x"82", -- 0x1F70
		x"2E",x"45",x"02",x"82",x"86",x"11",x"81",x"8C", -- 0x1F78
		x"31",x"12",x"4B",x"82",x"31",x"20",x"65",x"0F", -- 0x1F80
		x"44",x"A6",x"9B",x"40",x"65",x"C2",x"AC",x"36", -- 0x1F88
		x"0C",x"69",x"2E",x"A5",x"25",x"1F",x"81",x"74", -- 0x1F90
		x"14",x"46",x"F2",x"C3",x"29",x"55",x"BA",x"18", -- 0x1F98
		x"08",x"A5",x"22",x"75",x"C0",x"30",x"69",x"CA", -- 0x1FA0
		x"21",x"6A",x"AA",x"CF",x"60",x"FE",x"12",x"0C", -- 0x1FA8
		x"01",x"44",x"15",x"B0",x"86",x"EE",x"F2",x"19", -- 0x1FB0
		x"18",x"C3",x"10",x"B3",x"41",x"8C",x"22",x"40", -- 0x1FB8
		x"10",x"F9",x"5D",x"41",x"C4",x"00",x"6C",x"85", -- 0x1FC0
		x"69",x"00",x"42",x"35",x"DC",x"40",x"ED",x"20", -- 0x1FC8
		x"02",x"01",x"00",x"90",x"B2",x"39",x"9D",x"02", -- 0x1FD0
		x"50",x"62",x"12",x"38",x"EE",x"14",x"84",x"50", -- 0x1FD8
		x"C0",x"42",x"BE",x"4D",x"85",x"80",x"99",x"53", -- 0x1FE0
		x"2A",x"83",x"C1",x"D0",x"3F",x"51",x"5A",x"04", -- 0x1FE8
		x"89",x"DA",x"17",x"5E",x"8A",x"18",x"C0",x"10", -- 0x1FF0
		x"03",x"85",x"83",x"88",x"45",x"A7",x"05",x"01"  -- 0x1FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
