-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_L1 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_L1 is


	type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0000
		x"FE",x"FF",x"EF",x"FF",x"FE",x"EC",x"BC",x"F7", -- 0x0008
		x"CC",x"54",x"CD",x"FF",x"FE",x"FF",x"FF",x"FF", -- 0x0010
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0018
		x"DF",x"FF",x"FD",x"FF",x"AD",x"FF",x"A5",x"FF", -- 0x0020
		x"25",x"DD",x"8F",x"DD",x"78",x"D5",x"F8",x"FD", -- 0x0028
		x"00",x"73",x"00",x"FF",x"77",x"FF",x"A5",x"FF", -- 0x0030
		x"AD",x"FF",x"FD",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x0038
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0040
		x"DD",x"FF",x"EF",x"FF",x"FF",x"5C",x"CC",x"37", -- 0x0048
		x"CC",x"CC",x"DD",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x0050
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
		x"FF",x"FF",x"BB",x"FF",x"EF",x"FF",x"F7",x"FF", -- 0x0060
		x"77",x"FF",x"33",x"FF",x"80",x"3F",x"11",x"3D", -- 0x0068
		x"70",x"11",x"80",x"DD",x"91",x"DD",x"99",x"FF", -- 0x0070
		x"C8",x"FF",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0078
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0080
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DE",x"AF",x"E6", -- 0x0088
		x"CC",x"7E",x"CD",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x0090
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0098
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A0
		x"FF",x"DD",x"FF",x"DD",x"00",x"15",x"47",x"3D", -- 0x00A8
		x"77",x"BB",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00C0
		x"FF",x"FF",x"DD",x"FF",x"CC",x"DE",x"FF",x"FF", -- 0x00C8
		x"FF",x"EC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D8
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"8D",x"FF", -- 0x00E0
		x"88",x"DD",x"08",x"DD",x"77",x"DD",x"FF",x"FD", -- 0x00E8
		x"DD",x"33",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F0
		x"AB",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0100
		x"EF",x"FF",x"EF",x"FE",x"FF",x"6C",x"BB",x"FF", -- 0x0108
		x"CC",x"64",x"FF",x"FE",x"EF",x"FF",x"FF",x"FF", -- 0x0110
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0118
		x"DD",x"FF",x"AA",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x0120
		x"FF",x"DD",x"DD",x"DD",x"FF",x"5D",x"FF",x"FD", -- 0x0128
		x"00",x"73",x"DD",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x0130
		x"FF",x"FF",x"AA",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x0138
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0140
		x"FF",x"FF",x"FF",x"FF",x"FF",x"ED",x"FF",x"FF", -- 0x0148
		x"CC",x"DE",x"DD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0150
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0158
		x"DD",x"FF",x"AA",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0160
		x"77",x"DD",x"FF",x"DD",x"DD",x"95",x"FF",x"FD", -- 0x0168
		x"00",x"33",x"00",x"FF",x"88",x"FF",x"8D",x"FF", -- 0x0170
		x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0178
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0180
		x"DF",x"FF",x"CD",x"FF",x"CC",x"7E",x"9A",x"2E", -- 0x0188
		x"FF",x"CE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0190
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0198
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01A0
		x"FF",x"FF",x"F8",x"FF",x"11",x"BB",x"34",x"3D", -- 0x01A8
		x"08",x"91",x"FF",x"DD",x"FF",x"DD",x"FF",x"FF", -- 0x01B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01C0
		x"FD",x"FF",x"EF",x"FF",x"FF",x"4D",x"CC",x"BF", -- 0x01C8
		x"EF",x"EC",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x01E0
		x"AD",x"DD",x"AD",x"DD",x"F0",x"95",x"FF",x"FD", -- 0x01E8
		x"FF",x"33",x"87",x"FF",x"FC",x"FF",x"A9",x"FF", -- 0x01F0
		x"FB",x"FF",x"DD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0200
		x"FE",x"EE",x"EF",x"E6",x"EF",x"6F",x"ED",x"5E", -- 0x0208
		x"EE",x"64",x"EE",x"EE",x"EF",x"EE",x"FF",x"FF", -- 0x0210
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0218
		x"BB",x"FF",x"37",x"FF",x"FB",x"FF",x"FB",x"FF", -- 0x0220
		x"FB",x"FF",x"FB",x"FF",x"0E",x"FF",x"D4",x"77", -- 0x0228
		x"00",x"FF",x"33",x"FF",x"33",x"FF",x"77",x"FF", -- 0x0230
		x"73",x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"FF", -- 0x0238
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0240
		x"FF",x"FF",x"FF",x"DF",x"FF",x"CE",x"FF",x"65", -- 0x0248
		x"FF",x"CC",x"FF",x"DD",x"FF",x"FF",x"FF",x"FF", -- 0x0250
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0258
		x"FF",x"FF",x"BF",x"FF",x"FB",x"FF",x"FB",x"FF", -- 0x0260
		x"FB",x"FF",x"BF",x"FF",x"99",x"FF",x"51",x"FF", -- 0x0268
		x"11",x"FF",x"BB",x"FF",x"BB",x"FF",x"FB",x"FF", -- 0x0270
		x"FB",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0278
		x"FF",x"DD",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x0280
		x"FF",x"FF",x"FF",x"EE",x"EE",x"3F",x"DC",x"77", -- 0x0288
		x"EE",x"FF",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x0290
		x"FF",x"FF",x"FF",x"EE",x"FF",x"DD",x"FF",x"FF", -- 0x0298
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02A0
		x"77",x"77",x"66",x"77",x"AA",x"77",x"88",x"33", -- 0x02A8
		x"62",x"77",x"66",x"77",x"77",x"77",x"FF",x"FF", -- 0x02B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02B8
		x"FF",x"BB",x"FF",x"55",x"FF",x"FF",x"FF",x"EE", -- 0x02C0
		x"BB",x"FF",x"BB",x"BB",x"BB",x"FF",x"FB",x"FF", -- 0x02C8
		x"CC",x"00",x"FF",x"BB",x"FF",x"FF",x"FF",x"EE", -- 0x02D0
		x"FF",x"FF",x"FF",x"55",x"FF",x"BB",x"FF",x"FF", -- 0x02D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02E0
		x"FF",x"F7",x"F7",x"FF",x"62",x"FF",x"FF",x"FF", -- 0x02E8
		x"62",x"33",x"77",x"FF",x"F7",x"F7",x"FF",x"FF", -- 0x02F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02F8
		x"FF",x"BB",x"FF",x"9B",x"FF",x"99",x"FF",x"89", -- 0x0300
		x"FF",x"88",x"FF",x"88",x"EE",x"33",x"CC",x"11", -- 0x0308
		x"EE",x"00",x"FF",x"88",x"FF",x"88",x"FF",x"89", -- 0x0310
		x"FF",x"99",x"FF",x"9B",x"FF",x"BB",x"FF",x"FF", -- 0x0318
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0320
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"BF", -- 0x0328
		x"E6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0330
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0338
		x"FF",x"FF",x"FF",x"EF",x"FF",x"EF",x"FF",x"EF", -- 0x0340
		x"FF",x"EF",x"FF",x"EF",x"FF",x"FF",x"FF",x"EF", -- 0x0348
		x"FF",x"CC",x"FF",x"EE",x"FF",x"EE",x"FF",x"EF", -- 0x0350
		x"FF",x"EF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x0358
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0360
		x"BF",x"FF",x"FB",x"FF",x"FB",x"FF",x"5E",x"FF", -- 0x0368
		x"33",x"FF",x"FB",x"FF",x"BF",x"FF",x"FF",x"FF", -- 0x0370
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0378
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0380
		x"FF",x"7F",x"FF",x"F7",x"FF",x"A6",x"FE",x"3F", -- 0x0388
		x"FF",x"32",x"FF",x"77",x"FF",x"7F",x"FF",x"FF", -- 0x0390
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0398
		x"DD",x"FF",x"FF",x"FF",x"9F",x"FF",x"53",x"FF", -- 0x03A0
		x"DB",x"FF",x"DB",x"FF",x"3C",x"77",x"E2",x"B3", -- 0x03A8
		x"11",x"77",x"11",x"FF",x"77",x"FF",x"53",x"FF", -- 0x03B0
		x"9F",x"FF",x"FF",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x03B8
		x"FF",x"FF",x"CF",x"0F",x"CF",x"0F",x"CF",x"0F", -- 0x03C0
		x"CF",x"0F",x"CF",x"0F",x"CF",x"0F",x"CF",x"0F", -- 0x03C8
		x"EF",x"1F",x"CF",x"1F",x"CF",x"1F",x"CF",x"1F", -- 0x03D0
		x"CF",x"1F",x"EF",x"1F",x"FF",x"FF",x"FF",x"FF", -- 0x03D8
		x"FF",x"FF",x"0F",x"FF",x"0F",x"FF",x"0F",x"FF", -- 0x03E0
		x"0F",x"FF",x"0F",x"FF",x"0F",x"FF",x"0F",x"FF", -- 0x03E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03F8
		x"FF",x"FF",x"FF",x"10",x"FF",x"CD",x"FF",x"CD", -- 0x0400
		x"FF",x"98",x"BC",x"90",x"9A",x"90",x"FF",x"09", -- 0x0408
		x"FF",x"A9",x"FF",x"EF",x"FF",x"EF",x"FF",x"DC", -- 0x0410
		x"FF",x"94",x"FF",x"98",x"FF",x"FF",x"FF",x"FF", -- 0x0418
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"F7",x"FF", -- 0x0420
		x"D7",x"FF",x"B4",x"B7",x"B4",x"3B",x"4E",x"FF", -- 0x0428
		x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0430
		x"3D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0438
		x"FF",x"FF",x"FF",x"10",x"FF",x"FD",x"FF",x"FD", -- 0x0440
		x"CB",x"5D",x"FC",x"D5",x"DD",x"99",x"FF",x"91", -- 0x0448
		x"FF",x"FD",x"FF",x"DD",x"FF",x"EE",x"FF",x"FF", -- 0x0450
		x"FF",x"EE",x"FF",x"CC",x"FF",x"EE",x"FF",x"FF", -- 0x0458
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"77",x"FF", -- 0x0460
		x"D5",x"FF",x"E6",x"FF",x"D5",x"FF",x"33",x"FF", -- 0x0468
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0470
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0478
		x"FF",x"FF",x"FF",x"10",x"FF",x"DF",x"FF",x"DF", -- 0x0480
		x"FF",x"DD",x"FF",x"CC",x"FF",x"CC",x"FF",x"DD", -- 0x0488
		x"FF",x"DF",x"FF",x"CC",x"FF",x"FF",x"FF",x"FE", -- 0x0490
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"FF", -- 0x0498
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"F7",x"FF", -- 0x04A0
		x"F3",x"FF",x"F3",x"FF",x"F3",x"FF",x"7F",x"FF", -- 0x04A8
		x"77",x"FF",x"F7",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x04B0
		x"3D",x"FF",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04B8
		x"FF",x"FF",x"FF",x"10",x"FF",x"DD",x"FF",x"FF", -- 0x04C0
		x"EF",x"33",x"CE",x"33",x"EF",x"33",x"FF",x"3B", -- 0x04C8
		x"FF",x"DD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04D0
		x"FF",x"DD",x"FF",x"99",x"FF",x"FF",x"FF",x"FF", -- 0x04D8
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x04E0
		x"EE",x"FF",x"FF",x"77",x"66",x"FF",x"DD",x"FF", -- 0x04E8
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04F8
		x"FF",x"FF",x"FF",x"10",x"FF",x"DD",x"FF",x"DD", -- 0x0500
		x"9D",x"DD",x"FF",x"99",x"BB",x"DD",x"DD",x"DD", -- 0x0508
		x"FF",x"99",x"FF",x"DF",x"FF",x"FF",x"FF",x"DD", -- 0x0510
		x"FF",x"5D",x"FF",x"DD",x"FF",x"FF",x"FF",x"FF", -- 0x0518
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x0520
		x"FF",x"37",x"BB",x"FF",x"FF",x"BB",x"FF",x"77", -- 0x0528
		x"BB",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0530
		x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0538
		x"FF",x"FF",x"FF",x"10",x"FF",x"DD",x"FF",x"DD", -- 0x0540
		x"DD",x"FF",x"FF",x"DD",x"FF",x"FF",x"FF",x"FF", -- 0x0548
		x"FF",x"FF",x"FF",x"DD",x"FF",x"FF",x"FF",x"FF", -- 0x0550
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0558
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0560
		x"88",x"FF",x"88",x"77",x"88",x"FF",x"99",x"FF", -- 0x0568
		x"77",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0570
		x"77",x"FF",x"33",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0578
		x"FF",x"FF",x"FF",x"10",x"FF",x"CC",x"FF",x"EC", -- 0x0580
		x"FF",x"E8",x"FF",x"F8",x"FF",x"F8",x"FF",x"ED", -- 0x0588
		x"FF",x"CC",x"FF",x"EE",x"FF",x"FF",x"FF",x"CD", -- 0x0590
		x"FF",x"D4",x"FF",x"89",x"FF",x"FF",x"FF",x"FF", -- 0x0598
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"77",x"FF", -- 0x05A0
		x"7F",x"FF",x"77",x"FF",x"77",x"FF",x"77",x"FF", -- 0x05A8
		x"7F",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05B8
		x"FF",x"FF",x"FF",x"10",x"FF",x"DD",x"FF",x"DD", -- 0x05C0
		x"FF",x"75",x"EE",x"FD",x"FF",x"31",x"FF",x"99", -- 0x05C8
		x"FF",x"DD",x"FF",x"FF",x"FF",x"EF",x"FF",x"EE", -- 0x05D0
		x"FF",x"CC",x"FF",x"88",x"FF",x"EE",x"FF",x"FF", -- 0x05D8
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"7F",x"FF", -- 0x05E0
		x"34",x"7F",x"0F",x"7F",x"FF",x"77",x"33",x"FF", -- 0x05E8
		x"77",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F0
		x"77",x"FF",x"33",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x0600
		x"FF",x"DC",x"FF",x"CC",x"07",x"11",x"AA",x"10", -- 0x0608
		x"EE",x"01",x"FF",x"FD",x"FF",x"FF",x"FF",x"89", -- 0x0610
		x"FF",x"01",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x0618
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0620
		x"77",x"FF",x"7F",x"FF",x"8F",x"1D",x"FF",x"BB", -- 0x0628
		x"98",x"FF",x"77",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x0630
		x"11",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0640
		x"FF",x"FF",x"FF",x"DC",x"8E",x"10",x"FF",x"DC", -- 0x0648
		x"FF",x"DC",x"FF",x"99",x"FF",x"FF",x"FF",x"EE", -- 0x0650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0658
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0660
		x"FF",x"FF",x"F7",x"FF",x"87",x"3F",x"FF",x"FF", -- 0x0668
		x"F7",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"00", -- 0x0680
		x"FF",x"88",x"FF",x"EE",x"FF",x"CE",x"EF",x"55", -- 0x0688
		x"3B",x"99",x"FF",x"DD",x"FF",x"DD",x"FF",x"DF", -- 0x0690
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0698
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"11",x"FF", -- 0x06A0
		x"33",x"FF",x"FF",x"FF",x"77",x"FF",x"CD",x"FF", -- 0x06A8
		x"BB",x"9B",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x06B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"FF",x"5D", -- 0x06C0
		x"FF",x"DD",x"FF",x"FF",x"FF",x"FD",x"FF",x"D9", -- 0x06C8
		x"EE",x"DD",x"FF",x"DD",x"FF",x"99",x"FF",x"DD", -- 0x06D0
		x"FF",x"DD",x"FF",x"DD",x"FF",x"10",x"FF",x"FF", -- 0x06D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x06E0
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"BB",x"FF", -- 0x06E8
		x"EE",x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"FF", -- 0x06F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x0700
		x"FF",x"DD",x"FF",x"99",x"FF",x"FF",x"FF",x"DD", -- 0x0708
		x"FF",x"44",x"9D",x"00",x"00",x"00",x"FF",x"CC", -- 0x0710
		x"FF",x"CC",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x0718
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0720
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x0728
		x"DD",x"FF",x"99",x"37",x"00",x"11",x"77",x"FF", -- 0x0730
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0738
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x0740
		x"FF",x"FE",x"FF",x"EF",x"FF",x"59",x"FF",x"CC", -- 0x0748
		x"9F",x"00",x"FF",x"CC",x"FF",x"FF",x"FF",x"FF", -- 0x0750
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0758
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0760
		x"FF",x"FF",x"FF",x"FF",x"D3",x"FF",x"7F",x"FF", -- 0x0768
		x"47",x"3F",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x0780
		x"FF",x"ED",x"78",x"09",x"BB",x"10",x"FF",x"98", -- 0x0788
		x"FF",x"ED",x"FF",x"FE",x"FF",x"DD",x"FF",x"99", -- 0x0790
		x"FF",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A0
		x"77",x"FF",x"F8",x"D3",x"FF",x"BB",x"BB",x"FF", -- 0x07A8
		x"77",x"FF",x"FF",x"FF",x"F7",x"FF",x"3F",x"FF", -- 0x07B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B8
		x"FF",x"FF",x"EC",x"00",x"EC",x"00",x"FC",x"F0", -- 0x07C0
		x"EC",x"10",x"EC",x"D0",x"EC",x"10",x"FC",x"F0", -- 0x07C8
		x"FE",x"11",x"EC",x"71",x"FC",x"11",x"EC",x"71", -- 0x07D0
		x"FC",x"11",x"FE",x"F1",x"FF",x"FF",x"FF",x"FF", -- 0x07D8
		x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"60",x"FF", -- 0x07E0
		x"60",x"FF",x"00",x"FF",x"00",x"FF",x"F0",x"FF", -- 0x07E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F8
		x"FF",x"BF",x"FF",x"FB",x"FF",x"5B",x"FF",x"4A", -- 0x0800
		x"BB",x"5B",x"BB",x"BF",x"9A",x"F0",x"FB",x"F1", -- 0x0808
		x"EC",x"00",x"FF",x"00",x"FF",x"CC",x"FF",x"4A", -- 0x0810
		x"FF",x"5B",x"FF",x"FB",x"FF",x"BF",x"FF",x"FF", -- 0x0818
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0820
		x"FF",x"B7",x"FF",x"7B",x"7F",x"7B",x"EF",x"3D", -- 0x0828
		x"E6",x"33",x"FF",x"77",x"FF",x"B7",x"FF",x"FF", -- 0x0830
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0838
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"FF",x"55", -- 0x0840
		x"BB",x"EE",x"BB",x"FF",x"98",x"F0",x"FB",x"EF", -- 0x0848
		x"FC",x"00",x"FF",x"1F",x"FF",x"4A",x"FF",x"5B", -- 0x0850
		x"FF",x"FB",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF", -- 0x0858
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0860
		x"FF",x"FF",x"FF",x"FB",x"BB",x"BF",x"1D",x"FD", -- 0x0868
		x"62",x"33",x"FF",x"37",x"FF",x"FF",x"FF",x"FF", -- 0x0870
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0878
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0880
		x"BB",x"FF",x"BB",x"F1",x"9A",x"1F",x"FB",x"E9", -- 0x0888
		x"CF",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0890
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0898
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08A0
		x"FF",x"FB",x"FF",x"7F",x"67",x"FF",x"CF",x"95", -- 0x08A8
		x"7B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08B8
		x"FF",x"BB",x"FF",x"55",x"FF",x"FF",x"FF",x"FF", -- 0x08C0
		x"BB",x"EE",x"BB",x"FF",x"9A",x"BB",x"FB",x"FF", -- 0x08C8
		x"EC",x"00",x"FF",x"00",x"FF",x"11",x"FF",x"13", -- 0x08D0
		x"FF",x"37",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08E0
		x"FF",x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"FF", -- 0x08E8
		x"A6",x"33",x"FF",x"33",x"FF",x"FF",x"FF",x"FF", -- 0x08F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0900
		x"DF",x"FF",x"ED",x"FF",x"DC",x"7D",x"FC",x"0F", -- 0x0908
		x"ED",x"CE",x"DF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x0910
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0918
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x0920
		x"25",x"DD",x"AD",x"DD",x"F0",x"95",x"EF",x"7D", -- 0x0928
		x"00",x"73",x"FF",x"FF",x"AD",x"FF",x"25",x"FF", -- 0x0930
		x"AD",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0938
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"1B", -- 0x0940
		x"BB",x"01",x"BB",x"00",x"99",x"FF",x"FB",x"FF", -- 0x0948
		x"DD",x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x0950
		x"FF",x"FF",x"FF",x"55",x"FF",x"BB",x"FF",x"FF", -- 0x0958
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0960
		x"FF",x"FF",x"FF",x"BB",x"37",x"33",x"FF",x"FF", -- 0x0968
		x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0978
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0980
		x"BB",x"FF",x"BB",x"FF",x"A9",x"21",x"DA",x"79", -- 0x0988
		x"FC",x"80",x"FF",x"1F",x"FF",x"FF",x"FF",x"FF", -- 0x0990
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0998
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09A0
		x"FF",x"FF",x"FF",x"FF",x"B3",x"FF",x"2F",x"B5", -- 0x09A8
		x"E6",x"33",x"FF",x"37",x"FF",x"BF",x"FF",x"FF", -- 0x09B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"37",x"FF",x"17", -- 0x09C0
		x"BB",x"57",x"BB",x"47",x"88",x"67",x"EA",x"00", -- 0x09C8
		x"CC",x"E0",x"FF",x"00",x"FF",x"66",x"FF",x"55", -- 0x09D0
		x"FF",x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09E0
		x"FF",x"FB",x"FF",x"3F",x"67",x"BF",x"2E",x"57", -- 0x09E8
		x"66",x"33",x"FF",x"77",x"FF",x"BB",x"FF",x"FF", -- 0x09F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09F8
		x"FF",x"FF",x"FF",x"CE",x"FF",x"CF",x"FF",x"DE", -- 0x0A00
		x"FF",x"DE",x"FF",x"DE",x"FF",x"47",x"EE",x"B2", -- 0x0A08
		x"FF",x"00",x"FF",x"FC",x"FF",x"DD",x"FF",x"FE", -- 0x0A10
		x"FF",x"CF",x"FF",x"CE",x"FF",x"FF",x"FF",x"FF", -- 0x0A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A20
		x"77",x"77",x"6E",x"FF",x"7F",x"FF",x"F7",x"7B", -- 0x0A28
		x"A2",x"77",x"66",x"FF",x"77",x"77",x"FF",x"FF", -- 0x0A30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A38
		x"FF",x"FF",x"FF",x"DF",x"FF",x"DF",x"FF",x"DF", -- 0x0A40
		x"FF",x"DF",x"FF",x"DF",x"FF",x"9D",x"FF",x"A8", -- 0x0A48
		x"FF",x"88",x"FF",x"DD",x"FF",x"DD",x"FF",x"DF", -- 0x0A50
		x"FF",x"DF",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF", -- 0x0A58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A60
		x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"A6",x"FF", -- 0x0A68
		x"BB",x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"FF", -- 0x0A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x0A80
		x"EE",x"FF",x"EE",x"77",x"EE",x"55",x"CC",x"33", -- 0x0A88
		x"EE",x"44",x"EE",x"77",x"EE",x"EE",x"FF",x"FF", -- 0x0A90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A98
		x"BB",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AA0
		x"FF",x"FF",x"77",x"FF",x"EE",x"FF",x"DC",x"77", -- 0x0AA8
		x"00",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AB0
		x"FF",x"FF",x"77",x"FF",x"BB",x"FF",x"FF",x"FF", -- 0x0AB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AC0
		x"FF",x"FF",x"FF",x"FF",x"DD",x"FC",x"88",x"CE", -- 0x0AC8
		x"CC",x"EC",x"DD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AD8
		x"FF",x"FF",x"DC",x"FF",x"EA",x"FF",x"BB",x"FF", -- 0x0AE0
		x"B3",x"DD",x"33",x"DD",x"11",x"1D",x"E0",x"3D", -- 0x0AE8
		x"70",x"73",x"00",x"FF",x"88",x"FF",x"D8",x"FF", -- 0x0AF0
		x"FD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"FF", -- 0x0B08
		x"FF",x"23",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B18
		x"DD",x"FF",x"9D",x"FF",x"99",x"FF",x"99",x"FF", -- 0x0B20
		x"19",x"FF",x"11",x"FF",x"00",x"7F",x"00",x"37", -- 0x0B28
		x"F0",x"7F",x"11",x"FF",x"19",x"FF",x"99",x"FF", -- 0x0B30
		x"99",x"FF",x"9D",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x0B38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B40
		x"FF",x"FF",x"FF",x"DF",x"FF",x"DF",x"FF",x"0D", -- 0x0B48
		x"FF",x"CC",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF", -- 0x0B50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B58
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B60
		x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"7F",x"FF", -- 0x0B68
		x"3B",x"FF",x"77",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x0B70
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x0B78
		x"FF",x"FB",x"FF",x"B9",x"FF",x"BB",x"FF",x"BB", -- 0x0B80
		x"FF",x"AA",x"FF",x"BB",x"FF",x"77",x"EE",x"BC", -- 0x0B88
		x"FF",x"80",x"FF",x"88",x"FF",x"AA",x"FF",x"BB", -- 0x0B90
		x"FF",x"BB",x"FF",x"B9",x"FF",x"FB",x"FF",x"FF", -- 0x0B98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA0
		x"FE",x"FF",x"ED",x"FF",x"67",x"FF",x"FC",x"7F", -- 0x0BA8
		x"C4",x"FF",x"EC",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x0BB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB8
		x"FF",x"FF",x"DC",x"F0",x"DC",x"F0",x"CC",x"00", -- 0x0BC0
		x"DC",x"E0",x"DC",x"20",x"DC",x"E0",x"CC",x"00", -- 0x0BC8
		x"EE",x"F1",x"DC",x"91",x"CC",x"F1",x"DC",x"91", -- 0x0BD0
		x"CC",x"F1",x"EE",x"11",x"FF",x"FF",x"FF",x"FF", -- 0x0BD8
		x"FF",x"FF",x"F0",x"FF",x"F0",x"FF",x"90",x"FF", -- 0x0BE0
		x"90",x"FF",x"F0",x"FF",x"F0",x"FF",x"00",x"FF", -- 0x0BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF8
		x"FF",x"FF",x"FF",x"FE",x"FF",x"4D",x"FF",x"81", -- 0x0C00
		x"FF",x"CD",x"FF",x"EF",x"FF",x"DD",x"FF",x"B9", -- 0x0C08
		x"EE",x"99",x"EB",x"18",x"BC",x"18",x"EF",x"18", -- 0x0C10
		x"FF",x"DD",x"FF",x"FD",x"FF",x"10",x"FF",x"FF", -- 0x0C18
		x"FF",x"FF",x"FF",x"FF",x"D3",x"FF",x"FD",x"FF", -- 0x0C20
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"33",x"FF", -- 0x0C28
		x"6E",x"FF",x"87",x"FB",x"B4",x"B7",x"87",x"FF", -- 0x0C30
		x"F7",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C38
		x"FF",x"FF",x"FF",x"EF",x"FF",x"DD",x"FF",x"99", -- 0x0C40
		x"FF",x"DD",x"FF",x"EF",x"FF",x"EF",x"FF",x"ED", -- 0x0C48
		x"FF",x"C9",x"FF",x"A1",x"FE",x"21",x"FF",x"A1", -- 0x0C50
		x"FF",x"CD",x"FF",x"ED",x"FF",x"FE",x"FF",x"FF", -- 0x0C58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x0C68
		x"DD",x"FF",x"1F",x"77",x"FF",x"BB",x"00",x"77", -- 0x0C70
		x"7F",x"FF",x"F7",x"FF",x"11",x"FF",x"FF",x"FF", -- 0x0C78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"CD",x"FF",x"90", -- 0x0C80
		x"FF",x"CD",x"FF",x"FF",x"FF",x"EE",x"FF",x"DD", -- 0x0C88
		x"FF",x"DD",x"FF",x"9C",x"FF",x"9C",x"FF",x"8D", -- 0x0C90
		x"FF",x"DD",x"FF",x"DD",x"FF",x"10",x"FF",x"FF", -- 0x0C98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CA0
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"7F",x"FF", -- 0x0CA8
		x"7F",x"FF",x"77",x"FF",x"77",x"FF",x"77",x"FF", -- 0x0CB0
		x"7F",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"FF",x"DD", -- 0x0CC0
		x"FF",x"DD",x"FF",x"FF",x"FF",x"FD",x"FF",x"DD", -- 0x0CC8
		x"FF",x"77",x"EE",x"DD",x"DD",x"FF",x"EE",x"FF", -- 0x0CD0
		x"FF",x"DD",x"FF",x"DD",x"FF",x"10",x"FF",x"FF", -- 0x0CD8
		x"FF",x"FF",x"FF",x"FF",x"33",x"FF",x"77",x"FF", -- 0x0CE0
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x0CE8
		x"BB",x"FF",x"89",x"FF",x"88",x"7F",x"89",x"FF", -- 0x0CF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D00
		x"DF",x"FF",x"EF",x"FF",x"FF",x"5E",x"CC",x"26", -- 0x0D08
		x"CC",x"EC",x"FF",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x0D10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D18
		x"DD",x"FF",x"EA",x"FF",x"BB",x"FF",x"A3",x"FF", -- 0x0D20
		x"23",x"DD",x"33",x"DD",x"00",x"99",x"11",x"7D", -- 0x0D28
		x"07",x"73",x"80",x"FF",x"B3",x"FF",x"AA",x"FF", -- 0x0D30
		x"D8",x"FF",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"88",x"FF",x"CC", -- 0x0D40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"DD", -- 0x0D48
		x"FF",x"19",x"EF",x"11",x"EE",x"11",x"FF",x"11", -- 0x0D50
		x"FF",x"DD",x"FF",x"FD",x"FF",x"10",x"FF",x"FF", -- 0x0D58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FF", -- 0x0D60
		x"F7",x"FF",x"FF",x"FF",x"77",x"FF",x"BB",x"FF", -- 0x0D68
		x"EE",x"FF",x"BB",x"77",x"FF",x"BB",x"FF",x"77", -- 0x0D70
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D78
		x"FF",x"FF",x"FF",x"FE",x"FF",x"EF",x"FF",x"FE", -- 0x0D80
		x"FF",x"EE",x"FF",x"FF",x"FF",x"CE",x"FF",x"DF", -- 0x0D88
		x"FF",x"DF",x"FF",x"DC",x"FF",x"DC",x"FF",x"DC", -- 0x0D90
		x"FF",x"DF",x"FF",x"CC",x"FF",x"10",x"FF",x"FF", -- 0x0D98
		x"FF",x"FF",x"FF",x"FF",x"3D",x"FF",x"1D",x"FF", -- 0x0DA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FF", -- 0x0DA8
		x"FF",x"FF",x"7B",x"FF",x"7B",x"FF",x"7B",x"FF", -- 0x0DB0
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB8
		x"FF",x"FF",x"FF",x"FE",x"FF",x"EA",x"FF",x"CC", -- 0x0DC0
		x"FF",x"EE",x"FF",x"EF",x"FF",x"FD",x"FF",x"99", -- 0x0DC8
		x"FE",x"55",x"EF",x"5D",x"DE",x"D5",x"EF",x"5D", -- 0x0DD0
		x"FF",x"FD",x"FF",x"FD",x"FF",x"10",x"FF",x"FF", -- 0x0DD8
		x"FF",x"FF",x"FF",x"FF",x"13",x"FF",x"33",x"FF", -- 0x0DE0
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x0DE8
		x"3B",x"FF",x"D5",x"FF",x"E6",x"FF",x"E6",x"FF", -- 0x0DF0
		x"F7",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"45", -- 0x0E00
		x"FF",x"89",x"FF",x"EE",x"FF",x"DD",x"EE",x"98", -- 0x0E08
		x"47",x"98",x"BC",x"19",x"FF",x"CC",x"FF",x"DC", -- 0x0E10
		x"FF",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"FF", -- 0x0E20
		x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"6E",x"FF", -- 0x0E28
		x"4F",x"5D",x"7C",x"B7",x"FF",x"FF",x"77",x"FF", -- 0x0E30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E40
		x"FF",x"EE",x"FF",x"FF",x"FF",x"8D",x"FF",x"FE", -- 0x0E48
		x"FF",x"CC",x"78",x"10",x"FF",x"CE",x"FF",x"FF", -- 0x0E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E60
		x"FF",x"FF",x"FF",x"FF",x"3F",x"FF",x"FF",x"FF", -- 0x0E68
		x"FF",x"FF",x"34",x"D3",x"7F",x"FF",x"FF",x"FF", -- 0x0E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x0E80
		x"FF",x"DC",x"FF",x"CC",x"FF",x"DD",x"77",x"99", -- 0x0E88
		x"EE",x"DD",x"FF",x"CE",x"FF",x"EE",x"FF",x"88", -- 0x0E90
		x"FF",x"00",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x0E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EA0
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"DD", -- 0x0EA8
		x"EE",x"FF",x"77",x"FF",x"FF",x"FF",x"33",x"FF", -- 0x0EB0
		x"11",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EB8
		x"FF",x"FF",x"CC",x"00",x"CC",x"00",x"CC",x"00", -- 0x0EC0
		x"CC",x"00",x"CC",x"00",x"CC",x"00",x"CC",x"00", -- 0x0EC8
		x"EE",x"11",x"CC",x"11",x"CC",x"11",x"CC",x"11", -- 0x0ED0
		x"CC",x"11",x"EE",x"11",x"FF",x"FF",x"FF",x"FF", -- 0x0ED8
		x"FF",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"FF", -- 0x0EE0
		x"00",x"FF",x"00",x"FF",x"00",x"FF",x"00",x"FF", -- 0x0EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x0F00
		x"FF",x"CE",x"00",x"02",x"C8",x"02",x"FE",x"02", -- 0x0F08
		x"FF",x"DD",x"FF",x"FF",x"FF",x"99",x"FF",x"DD", -- 0x0F10
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F20
		x"77",x"FF",x"00",x"11",x"00",x"73",x"98",x"FF", -- 0x0F28
		x"F7",x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"FF", -- 0x0F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"CD",x"8F",x"8B", -- 0x0F48
		x"FF",x"DD",x"FF",x"49",x"FF",x"FE",x"FF",x"FE", -- 0x0F50
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F60
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"0F",x"3F", -- 0x0F68
		x"FF",x"FF",x"D3",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x0F80
		x"FF",x"89",x"FF",x"CD",x"FF",x"FF",x"FF",x"CD", -- 0x0F88
		x"FF",x"10",x"C9",x"18",x"77",x"01",x"FF",x"CD", -- 0x0F90
		x"FF",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA0
		x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x0FA8
		x"1D",x"FF",x"CF",x"73",x"FF",x"DD",x"77",x"FF", -- 0x0FB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB8
		x"FF",x"FF",x"DD",x"FF",x"DD",x"FF",x"CC",x"00", -- 0x0FC0
		x"DD",x"EE",x"DD",x"22",x"DD",x"EE",x"CC",x"00", -- 0x0FC8
		x"EE",x"FF",x"DD",x"99",x"CC",x"FF",x"DD",x"99", -- 0x0FD0
		x"CC",x"FF",x"EE",x"11",x"FF",x"FF",x"FF",x"FF", -- 0x0FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"99",x"FF", -- 0x0FE0
		x"99",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF", -- 0x0FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF8
		x"FF",x"EE",x"FF",x"DD",x"FF",x"CD",x"FF",x"CD", -- 0x1000
		x"FF",x"CD",x"FF",x"ED",x"FF",x"CD",x"DD",x"FF", -- 0x1008
		x"8A",x"CD",x"DF",x"02",x"EF",x"B3",x"ED",x"77", -- 0x1010
		x"EE",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1018
		x"FF",x"FF",x"77",x"FF",x"7F",x"FF",x"B3",x"FF", -- 0x1020
		x"E2",x"FF",x"7B",x"7B",x"7E",x"B3",x"E9",x"99", -- 0x1028
		x"81",x"55",x"12",x"7F",x"FC",x"F7",x"BA",x"B7", -- 0x1030
		x"EE",x"3F",x"FF",x"33",x"FF",x"FF",x"FF",x"FF", -- 0x1038
		x"FF",x"FF",x"FF",x"FF",x"FF",x"AD",x"FF",x"DE", -- 0x1040
		x"FF",x"8B",x"FF",x"EE",x"FF",x"CC",x"FF",x"FF", -- 0x1048
		x"FF",x"EF",x"CF",x"57",x"DD",x"73",x"EE",x"D5", -- 0x1050
		x"EF",x"9F",x"FF",x"9B",x"FF",x"FF",x"FF",x"FF", -- 0x1058
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"5D",x"F7", -- 0x1060
		x"BB",x"BB",x"74",x"D5",x"E9",x"FF",x"D2",x"F7", -- 0x1068
		x"96",x"F7",x"9A",x"D1",x"EE",x"9D",x"FF",x"FF", -- 0x1070
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1078
		x"FF",x"FF",x"FF",x"FF",x"DC",x"7F",x"CD",x"F3", -- 0x1080
		x"FF",x"C2",x"FF",x"2E",x"FF",x"CC",x"FF",x"DD", -- 0x1088
		x"FF",x"CD",x"FF",x"FF",x"EE",x"DF",x"CD",x"31", -- 0x1090
		x"EE",x"17",x"FF",x"72",x"FF",x"EE",x"FF",x"FF", -- 0x1098
		x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"24",x"77", -- 0x10A0
		x"42",x"BB",x"73",x"FF",x"E5",x"77",x"F0",x"F7", -- 0x10A8
		x"1E",x"B7",x"DD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10B0
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10C0
		x"DD",x"FF",x"FE",x"FF",x"FF",x"C5",x"CC",x"37", -- 0x10C8
		x"CC",x"5E",x"CD",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x10D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10D8
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"AD",x"FF", -- 0x10E0
		x"25",x"DD",x"E9",x"DD",x"F0",x"95",x"FF",x"B9", -- 0x10E8
		x"00",x"F3",x"77",x"FF",x"87",x"FF",x"AD",x"FF", -- 0x10F0
		x"AD",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10F8
		x"FF",x"FF",x"FF",x"EE",x"FF",x"C8",x"FF",x"BD", -- 0x1100
		x"FF",x"65",x"FF",x"BA",x"EE",x"D0",x"DE",x"85", -- 0x1108
		x"CF",x"0E",x"CC",x"11",x"FF",x"FF",x"FF",x"FF", -- 0x1110
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1118
		x"FF",x"FF",x"77",x"FF",x"DD",x"FF",x"34",x"77", -- 0x1120
		x"69",x"77",x"06",x"FF",x"3B",x"FF",x"B3",x"FF", -- 0x1128
		x"3B",x"FF",x"37",x"FF",x"99",x"77",x"A8",x"7F", -- 0x1130
		x"01",x"77",x"DC",x"FF",x"33",x"FF",x"FF",x"FF", -- 0x1138
		x"FF",x"FF",x"FF",x"BB",x"FF",x"77",x"FE",x"FE", -- 0x1140
		x"FF",x"DA",x"FE",x"61",x"FF",x"30",x"EF",x"98", -- 0x1148
		x"DE",x"08",x"ED",x"5D",x"DF",x"77",x"FF",x"FF", -- 0x1150
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1158
		x"FF",x"FF",x"99",x"FF",x"DB",x"FF",x"F3",x"FF", -- 0x1160
		x"D1",x"FF",x"3F",x"FF",x"3B",x"FF",x"F7",x"FF", -- 0x1168
		x"7F",x"FF",x"AE",x"3F",x"FD",x"3B",x"98",x"FF", -- 0x1170
		x"AE",x"7F",x"9D",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1178
		x"FF",x"FF",x"FF",x"FF",x"FF",x"66",x"EE",x"FF", -- 0x1180
		x"EE",x"54",x"FC",x"7C",x"DD",x"FA",x"EE",x"DE", -- 0x1188
		x"FF",x"00",x"EE",x"4C",x"EE",x"B7",x"DC",x"FF", -- 0x1190
		x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1198
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"F7",x"FF", -- 0x11A0
		x"B3",x"FF",x"3B",x"FF",x"3B",x"FF",x"7F",x"FF", -- 0x11A8
		x"FF",x"55",x"13",x"5D",x"DC",x"3B",x"CC",x"73", -- 0x11B0
		x"CD",x"77",x"CC",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"EF", -- 0x11D0
		x"7F",x"7F",x"7F",x"7F",x"1F",x"8F",x"1F",x"8F", -- 0x11D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x11F0
		x"BF",x"FF",x"BF",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x11F8
		x"FF",x"FF",x"FF",x"FF",x"CC",x"FF",x"DD",x"77", -- 0x1200
		x"DD",x"F5",x"FF",x"F3",x"EE",x"84",x"AA",x"10", -- 0x1208
		x"AA",x"61",x"CC",x"6F",x"ED",x"BC",x"FF",x"76", -- 0x1210
		x"FF",x"DC",x"FF",x"FF",x"FF",x"EE",x"FF",x"FF", -- 0x1218
		x"FF",x"FF",x"EE",x"FF",x"DD",x"77",x"CD",x"77", -- 0x1220
		x"EE",x"7B",x"DC",x"7F",x"8C",x"9D",x"3B",x"DD", -- 0x1228
		x"77",x"FF",x"7F",x"FF",x"3B",x"FF",x"BB",x"FF", -- 0x1230
		x"3B",x"FF",x"3B",x"FF",x"33",x"FF",x"73",x"FF", -- 0x1238
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1240
		x"FF",x"FF",x"AA",x"F7",x"9A",x"5D",x"DE",x"B6", -- 0x1248
		x"EF",x"B4",x"FF",x"79",x"AA",x"E2",x"DD",x"DD", -- 0x1250
		x"FE",x"AB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1258
		x"FF",x"FF",x"FF",x"FF",x"9D",x"FF",x"DF",x"7F", -- 0x1260
		x"BA",x"77",x"EC",x"BB",x"AE",x"3F",x"7F",x"FF", -- 0x1268
		x"FF",x"FF",x"33",x"FF",x"33",x"FF",x"1D",x"FF", -- 0x1270
		x"95",x"FF",x"5B",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1278
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1280
		x"FF",x"FF",x"FF",x"FF",x"AA",x"F7",x"ED",x"8C", -- 0x1288
		x"FA",x"80",x"EE",x"98",x"FF",x"13",x"DD",x"21", -- 0x1290
		x"EE",x"46",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF", -- 0x1298
		x"FF",x"FF",x"FF",x"FF",x"76",x"FF",x"9B",x"77", -- 0x12A0
		x"8D",x"7F",x"77",x"FF",x"BB",x"FF",x"7F",x"FF", -- 0x12A8
		x"FF",x"FF",x"95",x"FF",x"2E",x"FF",x"2C",x"FF", -- 0x12B0
		x"9A",x"77",x"EC",x"77",x"FF",x"FF",x"FF",x"FF", -- 0x12B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"EF", -- 0x12D0
		x"7F",x"FF",x"7F",x"BF",x"0F",x"0F",x"0F",x"4F", -- 0x12D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x12F0
		x"BF",x"FF",x"BF",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x12F8
		x"FF",x"FF",x"FF",x"EE",x"FF",x"C7",x"EE",x"2E", -- 0x1300
		x"EF",x"51",x"FF",x"99",x"FF",x"CE",x"FF",x"CD", -- 0x1308
		x"FF",x"89",x"FF",x"44",x"FF",x"CA",x"EE",x"E0", -- 0x1310
		x"CD",x"E2",x"CD",x"FF",x"FF",x"EE",x"FF",x"FF", -- 0x1318
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x1320
		x"FF",x"FF",x"FF",x"FF",x"EE",x"31",x"CF",x"95", -- 0x1328
		x"B4",x"7F",x"D6",x"77",x"B7",x"FF",x"AE",x"FF", -- 0x1330
		x"57",x"FF",x"31",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x1338
		x"FF",x"FF",x"FF",x"FF",x"FF",x"9B",x"EF",x"5F", -- 0x1340
		x"EE",x"95",x"CD",x"73",x"CF",x"57",x"FF",x"EF", -- 0x1348
		x"FF",x"EE",x"FF",x"CC",x"FF",x"CF",x"FF",x"9A", -- 0x1350
		x"FF",x"FC",x"FF",x"BD",x"FF",x"99",x"FF",x"FF", -- 0x1358
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1360
		x"FF",x"FF",x"EE",x"BF",x"BA",x"F3",x"D6",x"B7", -- 0x1368
		x"D3",x"7F",x"60",x"FF",x"30",x"77",x"19",x"FF", -- 0x1370
		x"5D",x"F7",x"EE",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x1378
		x"FF",x"FF",x"FF",x"FF",x"EE",x"77",x"EE",x"7F", -- 0x1380
		x"ED",x"FF",x"88",x"B3",x"FF",x"22",x"99",x"CD", -- 0x1388
		x"FF",x"CC",x"FF",x"DD",x"FF",x"CD",x"FF",x"CD", -- 0x1390
		x"FF",x"DC",x"FF",x"DC",x"FF",x"FF",x"FF",x"FF", -- 0x1398
		x"FF",x"FF",x"FF",x"FF",x"FF",x"33",x"EE",x"BF", -- 0x13A0
		x"FA",x"3B",x"74",x"7F",x"CF",x"77",x"B6",x"DD", -- 0x13A8
		x"69",x"99",x"11",x"3B",x"0C",x"FB",x"A2",x"FF", -- 0x13B0
		x"B3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13C8
		x"FF",x"FF",x"FF",x"FF",x"CF",x"0F",x"DF",x"FF", -- 0x13D0
		x"DF",x"FF",x"0F",x"0F",x"0F",x"0F",x"DF",x"FF", -- 0x13D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13E8
		x"FF",x"FF",x"FF",x"FF",x"3F",x"FF",x"BF",x"FF", -- 0x13F0
		x"BF",x"FF",x"3F",x"FF",x"3F",x"FF",x"FF",x"FF", -- 0x13F8
		x"FF",x"FF",x"FF",x"DD",x"FF",x"BD",x"EF",x"F0", -- 0x1400
		x"CC",x"BD",x"FF",x"35",x"FF",x"77",x"AB",x"F0", -- 0x1408
		x"47",x"0F",x"88",x"00",x"FF",x"00",x"FF",x"35", -- 0x1410
		x"CD",x"F0",x"CC",x"BD",x"FF",x"9F",x"FF",x"DD", -- 0x1418
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7D",x"FF", -- 0x1420
		x"BB",x"9D",x"77",x"FB",x"77",x"7B",x"BB",x"7F", -- 0x1428
		x"3E",x"D3",x"33",x"33",x"77",x"33",x"77",x"FB", -- 0x1430
		x"3B",x"9D",x"31",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1438
		x"FF",x"FF",x"FF",x"77",x"EF",x"CC",x"FF",x"C7", -- 0x1440
		x"DD",x"86",x"8B",x"D1",x"EE",x"5B",x"FF",x"34", -- 0x1448
		x"CD",x"A5",x"9A",x"48",x"9F",x"88",x"88",x"CC", -- 0x1450
		x"FF",x"BA",x"FF",x"9F",x"FF",x"88",x"FF",x"FF", -- 0x1458
		x"FF",x"FF",x"FF",x"FF",x"73",x"BB",x"EF",x"F7", -- 0x1460
		x"77",x"7F",x"EE",x"F3",x"32",x"33",x"84",x"77", -- 0x1468
		x"BB",x"DB",x"11",x"BB",x"22",x"FF",x"8E",x"F7", -- 0x1470
		x"95",x"FF",x"B3",x"FF",x"7F",x"FF",x"77",x"FF", -- 0x1478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"98", -- 0x1480
		x"DE",x"AC",x"CD",x"7B",x"EF",x"D1",x"DE",x"0C", -- 0x1488
		x"BB",x"AB",x"FF",x"47",x"EE",x"34",x"EE",x"AD", -- 0x1490
		x"FF",x"A6",x"EF",x"BB",x"FF",x"EE",x"FF",x"EE", -- 0x1498
		x"FF",x"FF",x"CD",x"77",x"EF",x"BB",x"CD",x"3B", -- 0x14A0
		x"FF",x"73",x"EE",x"C6",x"BA",x"9F",x"8E",x"BB", -- 0x14A8
		x"7B",x"CC",x"B7",x"FF",x"4C",x"FB",x"FB",x"7F", -- 0x14B0
		x"2D",x"B3",x"34",x"FF",x"2D",x"3B",x"AA",x"BB", -- 0x14B8
		x"FF",x"FF",x"FF",x"EE",x"FF",x"EE",x"FF",x"FF", -- 0x14C0
		x"FF",x"73",x"AA",x"7F",x"57",x"95",x"74",x"6E", -- 0x14C8
		x"BA",x"80",x"EF",x"99",x"B9",x"32",x"8A",x"BA", -- 0x14D0
		x"FF",x"8B",x"FF",x"57",x"FF",x"37",x"FF",x"33", -- 0x14D8
		x"FF",x"FF",x"3B",x"FF",x"DC",x"FF",x"98",x"BB", -- 0x14E0
		x"A9",x"7F",x"B9",x"7F",x"51",x"FF",x"77",x"FF", -- 0x14E8
		x"1D",x"B9",x"4A",x"9D",x"E1",x"F7",x"B4",x"B3", -- 0x14F0
		x"56",x"F3",x"BA",x"9F",x"DF",x"33",x"BB",x"FF", -- 0x14F8
		x"FF",x"77",x"FF",x"48",x"FF",x"CC",x"FF",x"FF", -- 0x1500
		x"FE",x"FF",x"EE",x"66",x"EE",x"08",x"FF",x"C4", -- 0x1508
		x"9A",x"C0",x"CF",x"84",x"FF",x"80",x"EE",x"6E", -- 0x1510
		x"EE",x"66",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x1518
		x"7F",x"77",x"F4",x"7F",x"97",x"FF",x"F7",x"FF", -- 0x1520
		x"FF",x"FB",x"3B",x"77",x"4C",x"BF",x"7B",x"FB", -- 0x1528
		x"F2",x"E0",x"E3",x"5B",x"C0",x"FB",x"3F",x"37", -- 0x1530
		x"7F",x"77",x"BB",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x1538
		x"FF",x"EE",x"FF",x"EF",x"EE",x"39",x"CD",x"18", -- 0x1540
		x"EE",x"98",x"FF",x"DD",x"FF",x"EE",x"FE",x"44", -- 0x1548
		x"EE",x"4C",x"EE",x"84",x"EE",x"EA",x"CC",x"CA", -- 0x1550
		x"DD",x"A4",x"DD",x"46",x"FF",x"AA",x"FF",x"FF", -- 0x1558
		x"BB",x"FF",x"3F",x"FF",x"3B",x"FF",x"76",x"FF", -- 0x1560
		x"EE",x"FF",x"66",x"7F",x"5D",x"6B",x"E3",x"5B", -- 0x1568
		x"5A",x"6A",x"61",x"AC",x"71",x"22",x"13",x"99", -- 0x1570
		x"8B",x"FF",x"89",x"FF",x"CC",x"FF",x"FF",x"FF", -- 0x1578
		x"FF",x"DD",x"FF",x"CE",x"FF",x"06",x"EE",x"97", -- 0x1580
		x"FF",x"51",x"DF",x"20",x"CC",x"45",x"FF",x"CC", -- 0x1588
		x"FF",x"EE",x"FF",x"95",x"FF",x"65",x"FF",x"9A", -- 0x1590
		x"FF",x"56",x"FF",x"46",x"FF",x"FF",x"FF",x"FF", -- 0x1598
		x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"CD",x"BB", -- 0x15A0
		x"FE",x"5F",x"45",x"A6",x"2F",x"D3",x"DA",x"1B", -- 0x15A8
		x"25",x"44",x"30",x"FF",x"89",x"F7",x"08",x"7F", -- 0x15B0
		x"EE",x"77",x"7F",x"FF",x"33",x"FF",x"FF",x"FF", -- 0x15B8
		x"FF",x"FF",x"DD",x"FE",x"FE",x"7F",x"EF",x"FF", -- 0x15C0
		x"FC",x"77",x"CC",x"C4",x"EE",x"12",x"BD",x"DD", -- 0x15C8
		x"DD",x"CC",x"FF",x"88",x"FF",x"97",x"FF",x"9A", -- 0x15D0
		x"FF",x"DC",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x15D8
		x"EE",x"FF",x"33",x"7F",x"BE",x"FF",x"16",x"BB", -- 0x15E0
		x"B8",x"1D",x"AD",x"77",x"E0",x"FF",x"5A",x"3B", -- 0x15E8
		x"21",x"95",x"11",x"9F",x"33",x"11",x"D5",x"FF", -- 0x15F0
		x"9F",x"FF",x"11",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EB",x"9B",x"DD", -- 0x1600
		x"FD",x"EE",x"ED",x"EE",x"EF",x"DD",x"BC",x"C7", -- 0x1608
		x"CC",x"CC",x"CC",x"EE",x"FD",x"EE",x"9B",x"CD", -- 0x1610
		x"FF",x"C8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1618
		x"BB",x"FF",x"DB",x"FF",x"F0",x"7F",x"DB",x"33", -- 0x1620
		x"CA",x"FF",x"EE",x"FF",x"F0",x"5D",x"0F",x"2E", -- 0x1628
		x"00",x"11",x"00",x"FF",x"CA",x"FF",x"F0",x"3B", -- 0x1630
		x"DB",x"33",x"9F",x"FF",x"BB",x"FF",x"FF",x"FF", -- 0x1638
		x"FF",x"EE",x"FF",x"CF",x"FF",x"DC",x"FF",x"9A", -- 0x1640
		x"FF",x"8F",x"FF",x"91",x"DD",x"CC",x"BD",x"89", -- 0x1648
		x"CE",x"9A",x"FE",x"C4",x"EC",x"77",x"EF",x"FF", -- 0x1650
		x"DC",x"7F",x"CC",x"77",x"FF",x"FF",x"FF",x"FF", -- 0x1658
		x"FF",x"FF",x"55",x"FF",x"9F",x"FF",x"95",x"FF", -- 0x1660
		x"E6",x"55",x"A9",x"1D",x"A5",x"99",x"7B",x"33", -- 0x1668
		x"88",x"FF",x"22",x"77",x"A9",x"95",x"DE",x"BB", -- 0x1670
		x"BE",x"3B",x"C4",x"3B",x"EE",x"33",x"FF",x"FF", -- 0x1678
		x"FF",x"DD",x"EE",x"D2",x"EE",x"79",x"FF",x"2D", -- 0x1680
		x"FE",x"7D",x"ED",x"03",x"FF",x"BA",x"FF",x"A9", -- 0x1688
		x"33",x"57",x"06",x"8C",x"37",x"B3",x"FE",x"77", -- 0x1690
		x"EC",x"3B",x"CD",x"7F",x"EE",x"3F",x"FF",x"FF", -- 0x1698
		x"3B",x"FF",x"BB",x"FF",x"66",x"3B",x"12",x"BB", -- 0x16A0
		x"5B",x"BB",x"F3",x"77",x"6E",x"FF",x"4C",x"77", -- 0x16A8
		x"03",x"B7",x"B8",x"7F",x"74",x"7F",x"CB",x"F7", -- 0x16B0
		x"D5",x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16B8
		x"FF",x"FF",x"FF",x"11",x"DD",x"37",x"CD",x"59", -- 0x16C0
		x"DD",x"E6",x"DD",x"84",x"CD",x"88",x"CD",x"11", -- 0x16C8
		x"FD",x"DD",x"FF",x"CD",x"FF",x"99",x"DD",x"A8", -- 0x16D0
		x"EF",x"73",x"DD",x"43",x"FF",x"77",x"FF",x"EE", -- 0x16D8
		x"FF",x"FF",x"BB",x"FF",x"17",x"FF",x"71",x"FF", -- 0x16E0
		x"9F",x"FF",x"62",x"55",x"A5",x"BF",x"78",x"D5", -- 0x16E8
		x"83",x"D5",x"99",x"0E",x"EF",x"88",x"DD",x"77", -- 0x16F0
		x"FD",x"FF",x"FF",x"FF",x"7F",x"FF",x"77",x"FF", -- 0x16F8
		x"FF",x"EE",x"FF",x"DD",x"CC",x"CD",x"CD",x"CD", -- 0x1700
		x"FE",x"10",x"9E",x"18",x"34",x"90",x"FE",x"89", -- 0x1708
		x"CD",x"01",x"CC",x"CD",x"FE",x"FF",x"FF",x"FE", -- 0x1710
		x"FF",x"98",x"EF",x"90",x"EE",x"EF",x"FF",x"FF", -- 0x1718
		x"FF",x"FF",x"77",x"FF",x"EE",x"FF",x"6E",x"7F", -- 0x1720
		x"91",x"F7",x"C7",x"B7",x"F4",x"D1",x"F7",x"F7", -- 0x1728
		x"99",x"7F",x"66",x"FF",x"FE",x"FF",x"FF",x"FF", -- 0x1730
		x"3F",x"FF",x"E9",x"FF",x"EE",x"FF",x"FF",x"FF", -- 0x1738
		x"FF",x"FF",x"FF",x"33",x"FF",x"37",x"FF",x"46", -- 0x1740
		x"FF",x"13",x"FF",x"B8",x"EC",x"98",x"BA",x"4D", -- 0x1748
		x"FE",x"48",x"8B",x"80",x"AA",x"F7",x"88",x"BB", -- 0x1750
		x"FF",x"FB",x"FF",x"FF",x"FF",x"EF",x"FF",x"EE", -- 0x1758
		x"FF",x"FF",x"BB",x"FF",x"FD",x"FF",x"A9",x"7F", -- 0x1760
		x"1E",x"7F",x"78",x"FF",x"E3",x"B3",x"84",x"7F", -- 0x1768
		x"3B",x"73",x"BB",x"FF",x"77",x"FF",x"D9",x"BB", -- 0x1770
		x"A9",x"7F",x"39",x"3B",x"19",x"FF",x"77",x"FF", -- 0x1778
		x"FF",x"FF",x"FF",x"EE",x"FF",x"66",x"DD",x"80", -- 0x1780
		x"DD",x"E3",x"EE",x"F9",x"EE",x"75",x"BB",x"23", -- 0x1788
		x"ED",x"11",x"BA",x"4C",x"DC",x"D1",x"AB",x"D5", -- 0x1790
		x"DF",x"15",x"BB",x"B9",x"FF",x"FF",x"FF",x"FF", -- 0x1798
		x"FF",x"FF",x"BB",x"FF",x"85",x"FF",x"78",x"FF", -- 0x17A0
		x"69",x"FF",x"D2",x"77",x"D5",x"FF",x"22",x"F7", -- 0x17A8
		x"FF",x"FF",x"BB",x"33",x"51",x"3F",x"B9",x"7F", -- 0x17B0
		x"98",x"FF",x"08",x"FF",x"15",x"FF",x"FF",x"FF", -- 0x17B8
		x"FF",x"FF",x"FF",x"9B",x"FF",x"CF",x"FF",x"BA", -- 0x17C0
		x"BB",x"23",x"8B",x"C3",x"99",x"78",x"CC",x"21", -- 0x17C8
		x"FF",x"00",x"FF",x"00",x"8B",x"95",x"DD",x"86", -- 0x17D0
		x"CD",x"E7",x"DD",x"CC",x"EE",x"77",x"FF",x"FF", -- 0x17D8
		x"BB",x"FF",x"7F",x"FF",x"B3",x"FF",x"95",x"FF", -- 0x17E0
		x"9F",x"FF",x"98",x"FF",x"33",x"BB",x"3B",x"53", -- 0x17E8
		x"8C",x"7F",x"32",x"F7",x"EE",x"73",x"EE",x"11", -- 0x17F0
		x"EF",x"3B",x"E7",x"77",x"FF",x"FF",x"FF",x"FF", -- 0x17F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"FF", -- 0x1800
		x"FF",x"CD",x"FF",x"FE",x"FF",x"CF",x"AB",x"F0", -- 0x1808
		x"47",x"C3",x"C8",x"00",x"FF",x"88",x"FF",x"FE", -- 0x1810
		x"FF",x"CD",x"FF",x"FF",x"FF",x"EE",x"FF",x"FF", -- 0x1818
		x"FF",x"FF",x"3D",x"FF",x"95",x"FF",x"95",x"FF", -- 0x1820
		x"95",x"FF",x"95",x"FF",x"1D",x"FF",x"E1",x"BB", -- 0x1828
		x"EF",x"F1",x"00",x"B3",x"00",x"FF",x"95",x"FF", -- 0x1830
		x"95",x"FF",x"95",x"FF",x"95",x"FF",x"3D",x"FF", -- 0x1838
		x"FF",x"91",x"FF",x"57",x"FF",x"42",x"FF",x"61", -- 0x1840
		x"FF",x"B4",x"FF",x"BC",x"FF",x"BC",x"FF",x"07", -- 0x1848
		x"EE",x"0F",x"CD",x"F3",x"8B",x"CC",x"FF",x"01", -- 0x1850
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1858
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1860
		x"77",x"FF",x"64",x"F7",x"AD",x"77",x"2E",x"FF", -- 0x1868
		x"DD",x"FF",x"33",x"FF",x"7B",x"FF",x"E0",x"FF", -- 0x1870
		x"79",x"FF",x"74",x"77",x"FF",x"77",x"FE",x"F7", -- 0x1878
		x"FF",x"FF",x"FF",x"77",x"EE",x"BB",x"FF",x"95", -- 0x1880
		x"EE",x"C2",x"FF",x"69",x"FF",x"E9",x"FF",x"24", -- 0x1888
		x"FF",x"CC",x"FF",x"01",x"FF",x"30",x"FF",x"61", -- 0x1890
		x"EE",x"0C",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x1898
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18A0
		x"CC",x"F7",x"10",x"FF",x"13",x"77",x"46",x"FF", -- 0x18A8
		x"4A",x"FF",x"A5",x"77",x"78",x"3B",x"BC",x"95", -- 0x18B0
		x"EF",x"F3",x"FF",x"77",x"FF",x"FF",x"FF",x"FF", -- 0x18B8
		x"FF",x"FF",x"FF",x"FF",x"CC",x"77",x"FE",x"BB", -- 0x18C0
		x"DC",x"E2",x"DD",x"4A",x"EE",x"1C",x"FF",x"CC", -- 0x18C8
		x"FF",x"30",x"FF",x"89",x"FF",x"F8",x"FF",x"02", -- 0x18D0
		x"FF",x"04",x"FF",x"DD",x"FF",x"BB",x"FF",x"FF", -- 0x18D8
		x"FF",x"FF",x"FF",x"FF",x"D8",x"FF",x"02",x"FF", -- 0x18E0
		x"F4",x"FF",x"73",x"FF",x"8E",x"FF",x"2D",x"BB", -- 0x18E8
		x"B4",x"A6",x"B4",x"D3",x"77",x"EE",x"77",x"FF", -- 0x18F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"FE", -- 0x1900
		x"FF",x"CC",x"C8",x"00",x"CF",x"0C",x"BC",x"C0", -- 0x1908
		x"EF",x"C0",x"FF",x"8C",x"FF",x"CC",x"FF",x"EE", -- 0x1910
		x"FF",x"EE",x"FF",x"EE",x"FF",x"FE",x"FF",x"FF", -- 0x1918
		x"FF",x"FF",x"F7",x"FF",x"F3",x"FF",x"B3",x"FF", -- 0x1920
		x"5D",x"FF",x"8C",x"10",x"CB",x"1F",x"5A",x"E1", -- 0x1928
		x"5A",x"B7",x"C3",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x1930
		x"3F",x"FF",x"7F",x"FF",x"BB",x"FF",x"77",x"FF", -- 0x1938
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"FF",x"51", -- 0x1940
		x"FF",x"E2",x"FF",x"A9",x"FF",x"89",x"FF",x"01", -- 0x1948
		x"DD",x"C0",x"FC",x"C0",x"47",x"68",x"88",x"00", -- 0x1950
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1958
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"91", -- 0x1960
		x"EC",x"48",x"47",x"B7",x"3C",x"F7",x"B4",x"BB", -- 0x1968
		x"B5",x"77",x"4A",x"FF",x"62",x"FF",x"60",x"FF", -- 0x1970
		x"13",x"FF",x"AB",x"FF",x"FD",x"FF",x"FF",x"FF", -- 0x1978
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"B3", -- 0x1980
		x"FF",x"40",x"FF",x"03",x"FF",x"99",x"FF",x"88", -- 0x1988
		x"FF",x"06",x"EE",x"78",x"CD",x"97",x"EF",x"5C", -- 0x1990
		x"DD",x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1998
		x"FF",x"FF",x"EE",x"FF",x"DC",x"3B",x"B8",x"BB", -- 0x19A0
		x"61",x"FF",x"69",x"77",x"3D",x"F7",x"5B",x"FF", -- 0x19A8
		x"35",x"F7",x"30",x"77",x"10",x"7F",x"CC",x"7F", -- 0x19B0
		x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"FF", -- 0x19C0
		x"EC",x"C1",x"CD",x"92",x"FE",x"07",x"FF",x"01", -- 0x19C8
		x"FF",x"00",x"FF",x"AC",x"EE",x"69",x"FF",x"D3", -- 0x19D0
		x"CD",x"D5",x"EC",x"BB",x"FF",x"FF",x"FF",x"FF", -- 0x19D8
		x"73",x"FF",x"FD",x"FF",x"D1",x"FF",x"D1",x"FF", -- 0x19E0
		x"D1",x"FF",x"D1",x"FF",x"1D",x"FF",x"E2",x"FF", -- 0x19E8
		x"B5",x"77",x"21",x"3B",x"A8",x"1D",x"76",x"77", -- 0x19F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19F8
		x"FF",x"8B",x"FF",x"9A",x"FF",x"9A",x"FF",x"9A", -- 0x1A00
		x"FF",x"9A",x"FF",x"8B",x"DD",x"78",x"BC",x"7F", -- 0x1A08
		x"DC",x"00",x"FF",x"00",x"FF",x"9A",x"FF",x"9A", -- 0x1A10
		x"FF",x"9A",x"FF",x"9A",x"FF",x"8B",x"FF",x"FF", -- 0x1A18
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"3B",x"FF", -- 0x1A20
		x"F7",x"FF",x"3F",x"FF",x"F0",x"5D",x"3C",x"2E", -- 0x1A28
		x"00",x"31",x"11",x"FF",x"F7",x"FF",x"3B",x"FF", -- 0x1A30
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A38
		x"FF",x"77",x"EE",x"FF",x"EE",x"E2",x"FF",x"E9", -- 0x1A40
		x"FF",x"70",x"FF",x"ED",x"FF",x"BB",x"FF",x"9A", -- 0x1A48
		x"FF",x"47",x"FF",x"59",x"DC",x"88",x"EC",x"E6", -- 0x1A50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"98", -- 0x1A60
		x"4C",x"8E",x"DE",x"3F",x"78",x"7F",x"1F",x"77", -- 0x1A68
		x"4C",x"FF",x"02",x"FF",x"E0",x"FF",x"68",x"FF", -- 0x1A70
		x"E8",x"FF",x"24",x"FF",x"EE",x"FF",x"98",x"FF", -- 0x1A78
		x"FF",x"FF",x"FF",x"FF",x"EA",x"FF",x"AD",x"5D", -- 0x1A80
		x"9A",x"D3",x"CD",x"C2",x"EE",x"0C",x"FF",x"01", -- 0x1A88
		x"FF",x"32",x"FF",x"07",x"EE",x"84",x"FE",x"FB", -- 0x1A90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A98
		x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"CD",x"7F", -- 0x1AA0
		x"21",x"77",x"71",x"FF",x"5A",x"FF",x"B7",x"FF", -- 0x1AA8
		x"4A",x"FF",x"79",x"FF",x"69",x"F7",x"34",x"FF", -- 0x1AB0
		x"9A",x"7F",x"CD",x"FB",x"EE",x"73",x"FF",x"FF", -- 0x1AB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AC0
		x"FF",x"EE",x"77",x"FE",x"BC",x"C0",x"56",x"A4", -- 0x1AC8
		x"DD",x"09",x"FF",x"51",x"FF",x"21",x"FF",x"97", -- 0x1AD0
		x"FF",x"62",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x1AD8
		x"FF",x"FF",x"DD",x"FF",x"AB",x"FF",x"02",x"FF", -- 0x1AE0
		x"34",x"FF",x"73",x"FF",x"7B",x"FF",x"E2",x"FF", -- 0x1AE8
		x"B5",x"FF",x"69",x"77",x"3C",x"BB",x"56",x"F7", -- 0x1AF0
		x"DD",x"7D",x"FF",x"FD",x"FF",x"F9",x"FF",x"FF", -- 0x1AF8
		x"FF",x"EE",x"FF",x"FD",x"FF",x"CD",x"FF",x"CD", -- 0x1B00
		x"FF",x"DC",x"FF",x"98",x"FF",x"18",x"DE",x"81", -- 0x1B08
		x"78",x"81",x"8F",x"19",x"80",x"11",x"FF",x"89", -- 0x1B10
		x"FF",x"FC",x"FF",x"DC",x"FF",x"EF",x"FF",x"FF", -- 0x1B18
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x1B20
		x"F7",x"FF",x"F7",x"FF",x"97",x"FF",x"B4",x"7F", -- 0x1B28
		x"B4",x"D3",x"87",x"3F",x"08",x"31",x"BB",x"FF", -- 0x1B30
		x"77",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B38
		x"FF",x"FF",x"FF",x"BB",x"FF",x"15",x"FF",x"A4", -- 0x1B40
		x"FF",x"F5",x"FF",x"70",x"FF",x"23",x"EE",x"49", -- 0x1B48
		x"CD",x"95",x"FE",x"A4",x"FC",x"4C",x"57",x"77", -- 0x1B50
		x"99",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B60
		x"99",x"B9",x"78",x"95",x"B4",x"39",x"B5",x"73", -- 0x1B68
		x"2E",x"FF",x"9D",x"FF",x"51",x"FF",x"F3",x"FF", -- 0x1B70
		x"B9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"77", -- 0x1B80
		x"CD",x"5D",x"EE",x"D3",x"EE",x"61",x"FF",x"12", -- 0x1B88
		x"FF",x"89",x"FE",x"8C",x"EE",x"4A",x"FD",x"C2", -- 0x1B90
		x"CD",x"95",x"FE",x"3B",x"EE",x"77",x"FF",x"FF", -- 0x1B98
		x"FF",x"FF",x"FF",x"FF",x"FE",x"F3",x"CC",x"BB", -- 0x1BA0
		x"67",x"B7",x"78",x"3B",x"E1",x"77",x"0E",x"FF", -- 0x1BA8
		x"95",x"FF",x"9D",x"FF",x"06",x"FF",x"31",x"FF", -- 0x1BB0
		x"98",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BC0
		x"AE",x"D5",x"D6",x"FE",x"C9",x"E1",x"DC",x"34", -- 0x1BC8
		x"FF",x"01",x"FF",x"20",x"FF",x"26",x"FF",x"61", -- 0x1BD0
		x"FF",x"71",x"FF",x"42",x"FF",x"37",x"FF",x"91", -- 0x1BD8
		x"FF",x"FF",x"FF",x"FF",x"AB",x"F7",x"65",x"FF", -- 0x1BE0
		x"79",x"FF",x"C2",x"FF",x"B7",x"FF",x"1D",x"FF", -- 0x1BE8
		x"BF",x"FF",x"42",x"FF",x"92",x"77",x"20",x"F7", -- 0x1BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF8
		x"FF",x"FF",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x1C00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"CF",x"0F", -- 0x1C08
		x"FF",x"99",x"FF",x"88",x"FF",x"88",x"FF",x"88", -- 0x1C10
		x"FF",x"88",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C18
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x1C20
		x"BB",x"FF",x"DF",x"77",x"FF",x"DD",x"0F",x"2E", -- 0x1C28
		x"3C",x"5D",x"33",x"FF",x"77",x"FF",x"77",x"FF", -- 0x1C30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C40
		x"FF",x"FF",x"FF",x"DD",x"EE",x"FF",x"BF",x"78", -- 0x1C48
		x"BF",x"10",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C60
		x"FF",x"FF",x"2E",x"FF",x"FF",x"DD",x"1F",x"EE", -- 0x1C68
		x"C0",x"31",x"52",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x1C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"98",x"FF",x"88", -- 0x1C80
		x"FF",x"88",x"FF",x"88",x"FF",x"EB",x"8F",x"7F", -- 0x1C88
		x"FF",x"88",x"FF",x"88",x"FF",x"FF",x"FF",x"FF", -- 0x1C90
		x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"FF",x"FF", -- 0x1C98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FF", -- 0x1CA0
		x"73",x"FF",x"31",x"FF",x"0F",x"5D",x"FF",x"EE", -- 0x1CA8
		x"12",x"31",x"30",x"7F",x"BB",x"FF",x"FF",x"FF", -- 0x1CB0
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CB8
		x"FF",x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CC0
		x"FF",x"FF",x"FF",x"77",x"DD",x"0F",x"8F",x"FF", -- 0x1CC8
		x"CC",x"80",x"FF",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1CD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"FF",x"FF", -- 0x1CD8
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x1CE0
		x"FF",x"FF",x"DD",x"FF",x"0F",x"5D",x"FF",x"EE", -- 0x1CE8
		x"00",x"31",x"11",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x1CF0
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF8
		x"FF",x"FF",x"FF",x"8B",x"FF",x"FF",x"FF",x"FF", -- 0x1D00
		x"FF",x"FF",x"9F",x"FF",x"8F",x"FF",x"8F",x"F8", -- 0x1D08
		x"FF",x"F8",x"FF",x"88",x"FF",x"88",x"FF",x"88", -- 0x1D10
		x"FF",x"C8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D18
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"7F",x"FF", -- 0x1D20
		x"BB",x"FF",x"BC",x"7F",x"FF",x"1D",x"B3",x"EE", -- 0x1D28
		x"00",x"31",x"11",x"FF",x"33",x"FF",x"77",x"FF", -- 0x1D30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D40
		x"BD",x"FF",x"9E",x"FE",x"8F",x"E3",x"FF",x"23", -- 0x1D48
		x"EE",x"00",x"FF",x"DC",x"FF",x"FF",x"FF",x"FF", -- 0x1D50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D60
		x"FF",x"FF",x"34",x"7F",x"0F",x"5D",x"F3",x"EE", -- 0x1D68
		x"40",x"31",x"10",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FF",x"8B", -- 0x1D80
		x"FF",x"8B",x"FF",x"8B",x"FF",x"8B",x"88",x"BF", -- 0x1D88
		x"FF",x"74",x"FF",x"FC",x"FF",x"FC",x"FF",x"FC", -- 0x1D90
		x"FF",x"FC",x"FF",x"8B",x"FF",x"FF",x"FF",x"FF", -- 0x1D98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DA0
		x"7F",x"FF",x"7F",x"FF",x"B4",x"5D",x"0F",x"2E", -- 0x1DA8
		x"D3",x"DD",x"84",x"F7",x"F7",x"FF",x"7F",x"FF", -- 0x1DB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"0F", -- 0x1DD0
		x"1F",x"0F",x"7F",x"7F",x"7F",x"7F",x"0F",x"0F", -- 0x1DD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x1DF0
		x"3F",x"FF",x"BF",x"FF",x"BF",x"FF",x"3F",x"FF", -- 0x1DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E00
		x"FF",x"FF",x"FF",x"EF",x"FF",x"EF",x"AB",x"D2", -- 0x1E08
		x"47",x"0F",x"BB",x"BC",x"FE",x"12",x"FF",x"FE", -- 0x1E10
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF", -- 0x1E20
		x"1D",x"FF",x"1D",x"FF",x"1D",x"FF",x"1D",x"FF", -- 0x1E28
		x"DF",x"11",x"E2",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x1E30
		x"F3",x"FF",x"F3",x"FF",x"1D",x"FF",x"FF",x"FF", -- 0x1E38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E40
		x"FF",x"FF",x"FF",x"FF",x"EF",x"D3",x"D9",x"0F", -- 0x1E48
		x"B3",x"DE",x"C8",x"40",x"FF",x"B0",x"FF",x"FF", -- 0x1E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E60
		x"FF",x"FF",x"FF",x"DB",x"F7",x"97",x"7E",x"1F", -- 0x1E68
		x"C2",x"FF",x"00",x"77",x"33",x"FF",x"FF",x"FF", -- 0x1E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x1E80
		x"FF",x"FF",x"FF",x"DD",x"EF",x"F3",x"AB",x"7F", -- 0x1E88
		x"77",x"98",x"C8",x"30",x"FF",x"88",x"FF",x"CC", -- 0x1E90
		x"FF",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E98
		x"FF",x"FF",x"FF",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x1EA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"9F",x"FF",x"1F", -- 0x1EA8
		x"F1",x"1F",x"D1",x"FF",x"11",x"FF",x"11",x"FF", -- 0x1EB0
		x"11",x"FF",x"31",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"FF", -- 0x1EC0
		x"FF",x"DD",x"FF",x"FF",x"FF",x"BB",x"AB",x"0F", -- 0x1EC8
		x"77",x"FF",x"C8",x"00",x"FF",x"88",x"FF",x"FF", -- 0x1ED0
		x"FF",x"DD",x"FF",x"FF",x"FF",x"EE",x"FF",x"FF", -- 0x1ED8
		x"FF",x"FF",x"DD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EE0
		x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"0F",x"BB", -- 0x1EE8
		x"FF",x"B9",x"00",x"73",x"00",x"FF",x"FF",x"FF", -- 0x1EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"FF", -- 0x1EF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F00
		x"FF",x"EE",x"FF",x"CC",x"FF",x"88",x"AB",x"0F", -- 0x1F08
		x"44",x"00",x"D9",x"FF",x"EF",x"F3",x"FF",x"DD", -- 0x1F10
		x"FF",x"FF",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x1F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"31",x"FF", -- 0x1F20
		x"11",x"FF",x"11",x"FF",x"51",x"FF",x"99",x"FF", -- 0x1F28
		x"00",x"11",x"FF",x"11",x"FF",x"99",x"FF",x"FF", -- 0x1F30
		x"FF",x"FF",x"FF",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x1F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"47",x"BB",x"FF", -- 0x1F48
		x"77",x"BC",x"C8",x"10",x"ED",x"D2",x"FF",x"FF", -- 0x1F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F60
		x"FF",x"FF",x"FF",x"FF",x"BB",x"FF",x"EE",x"F7", -- 0x1F68
		x"C2",x"FF",x"B1",x"1F",x"FF",x"9F",x"FF",x"DF", -- 0x1F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x1F80
		x"FF",x"FF",x"FF",x"DD",x"FE",x"77",x"BB",x"88", -- 0x1F88
		x"77",x"FF",x"C9",x"F1",x"FF",x"CC",x"FF",x"EE", -- 0x1F90
		x"FF",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F98
		x"FF",x"FF",x"FF",x"FF",x"55",x"FF",x"FF",x"FF", -- 0x1FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"33",x"FF", -- 0x1FA8
		x"EE",x"1F",x"51",x"17",x"11",x"9B",x"11",x"FF", -- 0x1FB0
		x"11",x"FF",x"11",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F", -- 0x1FD0
		x"7F",x"7F",x"7F",x"7F",x"0F",x"4F",x"0F",x"4F", -- 0x1FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"FF", -- 0x1FF0
		x"BF",x"FF",x"BF",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x1FF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2000
		x"06",x"FF",x"69",x"B7",x"F0",x"D3",x"F9",x"D3", -- 0x2008
		x"FF",x"DD",x"9F",x"3B",x"00",x"FF",x"FF",x"FF", -- 0x2010
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2018
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2020
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2028
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2030
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2038
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2040
		x"FF",x"FF",x"37",x"FF",x"E1",x"FF",x"78",x"7F", -- 0x2048
		x"8F",x"7F",x"00",x"FF",x"33",x"FF",x"FF",x"FF", -- 0x2050
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2058
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2060
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2068
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2070
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2078
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2080
		x"FF",x"FF",x"B1",x"FF",x"1F",x"FF",x"F4",x"7F", -- 0x2088
		x"11",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2090
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2098
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x20F8
		x"FF",x"33",x"EE",x"1D",x"FF",x"7B",x"CD",x"7B", -- 0x2100
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x2108
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x2110
		x"EF",x"6A",x"EF",x"5B",x"67",x"5B",x"EF",x"5B", -- 0x2118
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2120
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2128
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2130
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2138
		x"EF",x"5B",x"EF",x"5B",x"EF",x"5B",x"EF",x"4B", -- 0x2140
		x"EF",x"F0",x"EF",x"33",x"EF",x"48",x"EF",x"5B", -- 0x2148
		x"EF",x"5B",x"EF",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x2150
		x"EF",x"5B",x"0F",x"0F",x"F0",x"F0",x"0F",x"0F", -- 0x2158
		x"FF",x"DD",x"FF",x"DD",x"00",x"55",x"0F",x"DD", -- 0x2160
		x"F0",x"78",x"FF",x"77",x"00",x"77",x"77",x"FF", -- 0x2168
		x"77",x"FF",x"77",x"FF",x"77",x"FF",x"77",x"FF", -- 0x2170
		x"00",x"00",x"3C",x"87",x"F0",x"F0",x"1E",x"F3", -- 0x2178
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2180
		x"77",x"4A",x"EF",x"4A",x"EF",x"4A",x"EF",x"4A", -- 0x2188
		x"EF",x"4A",x"EF",x"4B",x"FE",x"F0",x"EF",x"33", -- 0x2190
		x"EF",x"48",x"EF",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x2198
		x"EF",x"3F",x"03",x"08",x"00",x"00",x"FF",x"FF", -- 0x21A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"FF",x"DD", -- 0x21A8
		x"00",x"55",x"0F",x"DD",x"F0",x"78",x"FF",x"77", -- 0x21B0
		x"00",x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x21B8
		x"67",x"7B",x"EF",x"7B",x"EF",x"6A",x"EF",x"7B", -- 0x21C0
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x21C8
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"CD",x"7B", -- 0x21D0
		x"FF",x"7B",x"EE",x"9D",x"FF",x"77",x"FF",x"FF", -- 0x21D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x21E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x21E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x21F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x21F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2200
		x"FF",x"FF",x"FF",x"77",x"FF",x"BF",x"FF",x"5B", -- 0x2208
		x"FF",x"5B",x"EF",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x2210
		x"CD",x"5B",x"EF",x"5B",x"EF",x"5B",x"EF",x"4A", -- 0x2218
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2220
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2228
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2230
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2238
		x"EF",x"5B",x"AB",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x2240
		x"EF",x"5B",x"EF",x"5B",x"67",x"4B",x"EF",x"F0", -- 0x2248
		x"EF",x"13",x"EF",x"48",x"EF",x"5B",x"EF",x"5B", -- 0x2250
		x"EF",x"5B",x"EF",x"0E",x"0F",x"0F",x"F0",x"F0", -- 0x2258
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2260
		x"FF",x"DD",x"00",x"DD",x"1F",x"55",x"C3",x"70", -- 0x2268
		x"FF",x"77",x"00",x"FF",x"77",x"FF",x"77",x"FF", -- 0x2270
		x"77",x"FF",x"00",x"00",x"3C",x"F0",x"F0",x"C3", -- 0x2278
		x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2280
		x"33",x"2E",x"67",x"5B",x"EF",x"5B",x"EF",x"4B", -- 0x2288
		x"EF",x"F0",x"67",x"33",x"EF",x"48",x"EF",x"4A", -- 0x2290
		x"EF",x"5B",x"EF",x"5B",x"AB",x"5B",x"EF",x"4A", -- 0x2298
		x"1E",x"B7",x"03",x"08",x"00",x"00",x"77",x"FF", -- 0x22A0
		x"77",x"FF",x"77",x"DD",x"00",x"DD",x"1F",x"55", -- 0x22A8
		x"E1",x"70",x"FF",x"77",x"00",x"FF",x"FF",x"FF", -- 0x22B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22B8
		x"EF",x"5B",x"EF",x"5B",x"EF",x"5B",x"CD",x"5B", -- 0x22C0
		x"EF",x"5B",x"EF",x"5B",x"EF",x"5B",x"FF",x"5B", -- 0x22C8
		x"FF",x"5B",x"FF",x"BF",x"FF",x"77",x"FF",x"FF", -- 0x22D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2300
		x"FF",x"FF",x"FF",x"77",x"FF",x"BF",x"FF",x"5B", -- 0x2308
		x"FF",x"5B",x"EF",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x2310
		x"CD",x"5B",x"EF",x"5B",x"EF",x"5B",x"EF",x"4A", -- 0x2318
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2320
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2328
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2330
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2338
		x"EF",x"5B",x"AB",x"5B",x"EF",x"5B",x"AF",x"5B", -- 0x2340
		x"EF",x"5B",x"CD",x"5B",x"67",x"4B",x"EF",x"F0", -- 0x2348
		x"AF",x"13",x"EF",x"48",x"EF",x"5B",x"6E",x"5B", -- 0x2350
		x"CF",x"5B",x"EF",x"0E",x"0E",x"0F",x"F0",x"B0", -- 0x2358
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2360
		x"FF",x"DD",x"00",x"DD",x"1F",x"55",x"C3",x"70", -- 0x2368
		x"FF",x"77",x"00",x"FF",x"77",x"FF",x"77",x"FF", -- 0x2370
		x"77",x"FF",x"00",x"00",x"3C",x"F0",x"F0",x"C3", -- 0x2378
		x"0F",x"0F",x"00",x"00",x"08",x"00",x"02",x"00", -- 0x2380
		x"11",x"2E",x"67",x"1B",x"AB",x"53",x"EF",x"4B", -- 0x2388
		x"CD",x"F0",x"EF",x"33",x"AE",x"48",x"EF",x"4A", -- 0x2390
		x"CD",x"5B",x"AA",x"5B",x"AB",x"5B",x"EF",x"4A", -- 0x2398
		x"1E",x"B7",x"03",x"08",x"00",x"00",x"77",x"FF", -- 0x23A0
		x"77",x"FF",x"77",x"DD",x"00",x"DD",x"1F",x"55", -- 0x23A8
		x"E1",x"70",x"FF",x"77",x"00",x"FF",x"FF",x"FF", -- 0x23B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23B8
		x"EF",x"5B",x"EF",x"5B",x"EF",x"5B",x"CD",x"5B", -- 0x23C0
		x"EF",x"5B",x"EF",x"5B",x"EF",x"5B",x"FF",x"5B", -- 0x23C8
		x"FF",x"5B",x"FF",x"BF",x"FF",x"77",x"FF",x"FF", -- 0x23D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2400
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2408
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2410
		x"FF",x"BC",x"FF",x"77",x"F0",x"F0",x"FF",x"FF", -- 0x2418
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x2420
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD", -- 0x2428
		x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"FF",x"77", -- 0x2430
		x"6E",x"FF",x"FF",x"0F",x"F0",x"F0",x"FF",x"C3", -- 0x2438
		x"FF",x"FF",x"FF",x"00",x"FF",x"8B",x"FF",x"FF", -- 0x2440
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2448
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2450
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2458
		x"FF",x"3F",x"00",x"06",x"66",x"00",x"FF",x"00", -- 0x2460
		x"FF",x"88",x"FF",x"88",x"FF",x"DD",x"FF",x"DD", -- 0x2468
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x2470
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2480
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2488
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x2490
		x"BB",x"FF",x"BB",x"DE",x"BB",x"BB",x"E1",x"0F", -- 0x2498
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24A8
		x"FF",x"FF",x"FF",x"EE",x"FF",x"FF",x"FF",x"DD", -- 0x24B0
		x"FF",x"BB",x"7F",x"77",x"FF",x"3C",x"0F",x"3C", -- 0x24B8
		x"00",x"FF",x"33",x"88",x"33",x"CD",x"BB",x"FF", -- 0x24C0
		x"BB",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x24C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24D8
		x"FF",x"8F",x"00",x"03",x"77",x"00",x"FF",x"88", -- 0x24E0
		x"FF",x"CC",x"FF",x"EE",x"FF",x"EE",x"FF",x"FF", -- 0x24E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2500
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2508
		x"FF",x"FF",x"FF",x"EE",x"FF",x"DD",x"FF",x"EF", -- 0x2510
		x"FF",x"EF",x"FF",x"AB",x"FF",x"EF",x"FF",x"EF", -- 0x2518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2520
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2528
		x"FF",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x2530
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2538
		x"FF",x"EF",x"FF",x"EF",x"FF",x"67",x"FF",x"27", -- 0x2540
		x"FF",x"67",x"FF",x"67",x"FF",x"47",x"EE",x"03", -- 0x2548
		x"EE",x"6E",x"FF",x"EF",x"FF",x"67",x"EE",x"67", -- 0x2550
		x"EE",x"67",x"01",x"23",x"1E",x"C1",x"CF",x"0F", -- 0x2558
		x"BB",x"FF",x"BB",x"FF",x"BB",x"FF",x"BB",x"FF", -- 0x2560
		x"BB",x"DD",x"BB",x"DD",x"88",x"DD",x"0F",x"70", -- 0x2568
		x"EE",x"77",x"00",x"FF",x"99",x"FF",x"99",x"FF", -- 0x2570
		x"99",x"FF",x"88",x"00",x"F0",x"C3",x"07",x"D3", -- 0x2578
		x"01",x"01",x"08",x"00",x"9B",x"00",x"FF",x"33", -- 0x2580
		x"FF",x"67",x"EE",x"CF",x"EE",x"23",x"EE",x"47", -- 0x2588
		x"FF",x"6E",x"FF",x"67",x"FF",x"45",x"FF",x"27", -- 0x2590
		x"FF",x"67",x"FF",x"EF",x"FF",x"EF",x"FF",x"EF", -- 0x2598
		x"01",x"0C",x"00",x"00",x"11",x"FF",x"11",x"FF", -- 0x25A0
		x"99",x"DD",x"DD",x"DD",x"CC",x"55",x"0F",x"70", -- 0x25A8
		x"EE",x"77",x"00",x"FF",x"BB",x"FF",x"BB",x"FF", -- 0x25B0
		x"BB",x"FF",x"BB",x"FF",x"BB",x"FF",x"FF",x"FF", -- 0x25B8
		x"FF",x"EF",x"FF",x"AB",x"FF",x"EF",x"FF",x"EF", -- 0x25C0
		x"FF",x"DD",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x25C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25E0
		x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2600
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2608
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2610
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x2618
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2620
		x"FF",x"FF",x"EE",x"FF",x"DD",x"3B",x"DD",x"7F", -- 0x2628
		x"DD",x"5D",x"DD",x"5D",x"DD",x"5D",x"DD",x"5D", -- 0x2630
		x"DD",x"4C",x"DD",x"4C",x"59",x"0F",x"E3",x"F0", -- 0x2638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2640
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2658
		x"0C",x"00",x"CC",x"00",x"CC",x"00",x"CC",x"55", -- 0x2660
		x"CC",x"5D",x"DD",x"5D",x"DD",x"5D",x"DD",x"7F", -- 0x2668
		x"DD",x"3B",x"EE",x"77",x"FF",x"FF",x"FF",x"FF", -- 0x2670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2680
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2688
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2690
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2698
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26A8
		x"FF",x"FF",x"FF",x"AB",x"FF",x"AB",x"FF",x"AB", -- 0x26B0
		x"FF",x"AB",x"FF",x"AB",x"FF",x"AB",x"EF",x"D6", -- 0x26B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26D8
		x"EF",x"08",x"FF",x"88",x"FF",x"88",x"FF",x"89", -- 0x26E0
		x"FF",x"AB",x"FF",x"AB",x"FF",x"AB",x"FF",x"FF", -- 0x26E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2700
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2708
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x2710
		x"BB",x"FF",x"BB",x"DE",x"BB",x"BB",x"E1",x"0F", -- 0x2718
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2720
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2728
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF", -- 0x2730
		x"FF",x"BB",x"7F",x"57",x"BB",x"3C",x"0F",x"3C", -- 0x2738
		x"00",x"FF",x"33",x"88",x"33",x"CD",x"BB",x"FF", -- 0x2740
		x"BB",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x2748
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2750
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2758
		x"FF",x"8F",x"02",x"03",x"77",x"00",x"FF",x"BF", -- 0x2760
		x"FF",x"EE",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x2768
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2788
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2790
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27A8
		x"FF",x"FF",x"FF",x"AB",x"FF",x"AB",x"FF",x"CD", -- 0x27B0
		x"FF",x"EF",x"FF",x"8B",x"FF",x"AF",x"EF",x"D6", -- 0x27B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27D8
		x"EF",x"08",x"FF",x"89",x"FF",x"CC",x"FF",x"8C", -- 0x27E0
		x"FF",x"AB",x"FF",x"8B",x"FF",x"AB",x"FF",x"FF", -- 0x27E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2800
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2808
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2810
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2818
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2820
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2828
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2830
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2838
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2840
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2848
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2850
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2858
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2860
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2868
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2870
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2878
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2880
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2888
		x"FF",x"FF",x"FF",x"FF",x"FF",x"15",x"FF",x"37", -- 0x2890
		x"FF",x"AE",x"FF",x"2A",x"FE",x"26",x"DE",x"78", -- 0x2898
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28B0
		x"FF",x"FF",x"EF",x"E6",x"DD",x"CF",x"F3",x"FF", -- 0x28B8
		x"EF",x"02",x"FF",x"08",x"FF",x"22",x"FF",x"37", -- 0x28C0
		x"FF",x"15",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28D8
		x"CC",x"00",x"EE",x"6E",x"FF",x"FF",x"FF",x"FF", -- 0x28E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2900
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2908
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"BB", -- 0x2910
		x"FF",x"DF",x"FF",x"57",x"FF",x"DF",x"FF",x"CE", -- 0x2918
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2920
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2928
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2930
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2938
		x"FF",x"DF",x"FF",x"DF",x"FE",x"DF",x"EE",x"DF", -- 0x2940
		x"EE",x"57",x"EE",x"DF",x"EE",x"DF",x"EC",x"DF", -- 0x2948
		x"CC",x"89",x"CC",x"E8",x"CC",x"98",x"C8",x"46", -- 0x2950
		x"CC",x"DF",x"88",x"DF",x"00",x"00",x"78",x"70", -- 0x2958
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2960
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"FF", -- 0x2968
		x"7C",x"F7",x"22",x"FF",x"E2",x"FF",x"66",x"FF", -- 0x2970
		x"77",x"FF",x"77",x"FF",x"FF",x"DD",x"C3",x"7A", -- 0x2978
		x"07",x"0B",x"B0",x"F0",x"88",x"00",x"CC",x"FF", -- 0x2980
		x"CC",x"57",x"EE",x"99",x"EC",x"AB",x"CC",x"40", -- 0x2988
		x"EC",x"CC",x"EE",x"DF",x"EE",x"57",x"EE",x"DF", -- 0x2990
		x"EE",x"57",x"FE",x"9B",x"FF",x"DF",x"FF",x"DF", -- 0x2998
		x"F3",x"CD",x"F0",x"95",x"77",x"FF",x"77",x"FF", -- 0x29A0
		x"77",x"FF",x"BB",x"FF",x"7F",x"FF",x"30",x"F7", -- 0x29A8
		x"E2",x"FF",x"EE",x"FF",x"EE",x"FF",x"FF",x"FF", -- 0x29B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29B8
		x"FF",x"CE",x"FF",x"DF",x"FF",x"57",x"FF",x"DF", -- 0x29C0
		x"FF",x"BB",x"FF",x"D9",x"FF",x"FF",x"FF",x"FF", -- 0x29C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"FF",x"FE", -- 0x2A10
		x"FF",x"CC",x"FF",x"AA",x"FF",x"CC",x"FF",x"A4", -- 0x2A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A30
		x"FF",x"FF",x"FF",x"BD",x"F6",x"00",x"3F",x"8D", -- 0x2A38
		x"FF",x"4F",x"FF",x"88",x"FF",x"88",x"FF",x"AA", -- 0x2A40
		x"FF",x"98",x"FF",x"DD",x"FF",x"FF",x"FF",x"FF", -- 0x2A48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A58
		x"CC",x"77",x"76",x"F0",x"FF",x"9F",x"FF",x"FF", -- 0x2A60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"EC", -- 0x2A90
		x"FF",x"EE",x"FF",x"EF",x"FF",x"CC",x"FF",x"DA", -- 0x2A98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FF", -- 0x2AB0
		x"77",x"FF",x"77",x"FD",x"73",x"55",x"17",x"EE", -- 0x2AB8
		x"FF",x"CC",x"FF",x"CC",x"FF",x"FF",x"FF",x"EC", -- 0x2AC0
		x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AD8
		x"33",x"80",x"FF",x"DF",x"FF",x"FF",x"F7",x"FF", -- 0x2AE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B10
		x"FF",x"D9",x"FF",x"BB",x"FF",x"BB",x"FF",x"F7", -- 0x2B18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B38
		x"FF",x"76",x"FF",x"66",x"FF",x"66",x"FF",x"22", -- 0x2B40
		x"FF",x"66",x"FF",x"66",x"FE",x"66",x"EE",x"00", -- 0x2B48
		x"EE",x"66",x"EE",x"45",x"EE",x"66",x"EC",x"66", -- 0x2B50
		x"CC",x"22",x"88",x"22",x"DD",x"FF",x"07",x"03", -- 0x2B58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B68
		x"BB",x"FF",x"7C",x"FF",x"91",x"FF",x"55",x"FF", -- 0x2B70
		x"F7",x"FF",x"F7",x"FF",x"FE",x"77",x"F7",x"FB", -- 0x2B78
		x"00",x"00",x"88",x"00",x"CC",x"66",x"EC",x"22", -- 0x2B80
		x"EE",x"66",x"EE",x"45",x"FE",x"10",x"FF",x"66", -- 0x2B88
		x"FF",x"66",x"FF",x"22",x"FF",x"66",x"FF",x"66", -- 0x2B90
		x"FF",x"66",x"FF",x"76",x"FF",x"B3",x"FF",x"BB", -- 0x2B98
		x"01",x"F7",x"77",x"FF",x"77",x"FF",x"F7",x"FF", -- 0x2BA0
		x"BB",x"FF",x"7C",x"FF",x"91",x"FF",x"DD",x"FF", -- 0x2BA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BB8
		x"FF",x"BB",x"FF",x"BB",x"FF",x"D9",x"FF",x"FF", -- 0x2BC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"FF", -- 0x2CB0
		x"AA",x"FF",x"DD",x"FF",x"DD",x"EC",x"4F",x"99", -- 0x2CB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CD8
		x"88",x"FC",x"FD",x"FF",x"88",x"FF",x"DD",x"FF", -- 0x2CE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD", -- 0x2D18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D38
		x"FF",x"FD",x"FF",x"DC",x"FF",x"EA",x"FF",x"AA", -- 0x2D40
		x"FF",x"AA",x"FF",x"AA",x"FF",x"AA",x"FF",x"80", -- 0x2D48
		x"FF",x"22",x"FF",x"22",x"FE",x"51",x"EE",x"22", -- 0x2D50
		x"EE",x"00",x"FC",x"A2",x"00",x"00",x"37",x"BB", -- 0x2D58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D68
		x"FF",x"FF",x"73",x"FF",x"7C",x"FF",x"91",x"FF", -- 0x2D70
		x"55",x"FF",x"F7",x"FF",x"10",x"FF",x"F7",x"F7", -- 0x2D78
		x"E0",x"F0",x"CC",x"00",x"EE",x"80",x"FE",x"33", -- 0x2D80
		x"FE",x"23",x"FF",x"10",x"FF",x"22",x"FF",x"80", -- 0x2D88
		x"FF",x"AA",x"FF",x"AA",x"FF",x"AA",x"FF",x"AA", -- 0x2D90
		x"FF",x"EA",x"FF",x"DC",x"FF",x"FD",x"FF",x"FF", -- 0x2D98
		x"E0",x"FF",x"77",x"FF",x"F7",x"FF",x"73",x"FF", -- 0x2DA0
		x"7C",x"FF",x"91",x"FF",x"DD",x"FF",x"FF",x"FF", -- 0x2DA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DF8
		x"FF",x"B9",x"FF",x"D5",x"FF",x"15",x"FF",x"9D", -- 0x2E00
		x"FF",x"9D",x"FE",x"9D",x"EE",x"9D",x"FF",x"9D", -- 0x2E08
		x"FF",x"9D",x"FF",x"BF",x"FD",x"8F",x"DD",x"8C", -- 0x2E10
		x"D9",x"9D",x"91",x"8C",x"FF",x"F9",x"7C",x"F0", -- 0x2E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E28
		x"FF",x"FF",x"BB",x"FF",x"7D",x"FF",x"51",x"FF", -- 0x2E30
		x"DD",x"FF",x"DD",x"FF",x"EE",x"FF",x"97",x"F7", -- 0x2E38
		x"00",x"06",x"F0",x"F0",x"F8",x"75",x"FD",x"9D", -- 0x2E40
		x"FD",x"8F",x"FF",x"8C",x"FF",x"9D",x"FF",x"9D", -- 0x2E48
		x"EE",x"9D",x"FE",x"9D",x"FF",x"9D",x"FF",x"9D", -- 0x2E50
		x"FF",x"15",x"FF",x"D5",x"FF",x"B9",x"FF",x"FF", -- 0x2E58
		x"10",x"77",x"FF",x"77",x"FF",x"77",x"BB",x"FF", -- 0x2E60
		x"7D",x"FF",x"51",x"FF",x"DD",x"FF",x"DD",x"FF", -- 0x2E68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E88
		x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"EE", -- 0x2E90
		x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EA8
		x"FF",x"FF",x"B7",x"FF",x"73",x"FF",x"F7",x"FF", -- 0x2EB0
		x"FF",x"FF",x"7F",x"FF",x"5F",x"B3",x"FF",x"CF", -- 0x2EB8
		x"FF",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC0
		x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x2EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED8
		x"11",x"80",x"BB",x"FF",x"7F",x"FF",x"7F",x"FF", -- 0x2EE0
		x"FF",x"FF",x"B7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF8
		x"FF",x"33",x"FE",x"FD",x"EE",x"5D",x"FF",x"5D", -- 0x2F00
		x"FF",x"5D",x"FD",x"5D",x"DD",x"5D",x"DD",x"5D", -- 0x2F08
		x"DD",x"5D",x"D9",x"5D",x"99",x"5D",x"91",x"5D", -- 0x2F10
		x"91",x"5D",x"77",x"FF",x"87",x"C3",x"F0",x"E1", -- 0x2F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F30
		x"FF",x"FF",x"44",x"FF",x"8B",x"FF",x"BB",x"F3", -- 0x2F38
		x"08",x"0C",x"F0",x"F0",x"F0",x"F1",x"F1",x"FD", -- 0x2F40
		x"99",x"5D",x"D9",x"5D",x"DD",x"5D",x"DD",x"5D", -- 0x2F48
		x"DD",x"5D",x"FD",x"5D",x"FF",x"5D",x"FF",x"5D", -- 0x2F50
		x"EE",x"5D",x"FE",x"FD",x"FF",x"33",x"FF",x"FF", -- 0x2F58
		x"40",x"77",x"F4",x"77",x"FF",x"77",x"FF",x"77", -- 0x2F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F88
		x"FF",x"FF",x"FF",x"B3",x"FF",x"55",x"FF",x"66", -- 0x2F90
		x"FF",x"57",x"FF",x"57",x"FF",x"DF",x"FF",x"AD", -- 0x2F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FB0
		x"FF",x"FE",x"77",x"EC",x"EC",x"8F",x"7F",x"FE", -- 0x2FB8
		x"FF",x"98",x"FF",x"31",x"FF",x"53",x"FF",x"C6", -- 0x2FC0
		x"FF",x"55",x"FF",x"B3",x"FF",x"FF",x"FF",x"FF", -- 0x2FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD8
		x"EC",x"00",x"77",x"FC",x"FF",x"FE",x"FF",x"FF", -- 0x2FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FF8
		x"FF",x"33",x"EE",x"1D",x"FF",x"7B",x"CD",x"7B", -- 0x3000
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3008
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3010
		x"EF",x"6A",x"EF",x"5B",x"67",x"5B",x"EF",x"5B", -- 0x3018
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3020
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3028
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3030
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3038
		x"EF",x"5B",x"EF",x"5B",x"EF",x"5B",x"EF",x"4B", -- 0x3040
		x"EF",x"B4",x"EF",x"37",x"EF",x"48",x"ED",x"1B", -- 0x3048
		x"FE",x"5A",x"EF",x"A1",x"68",x"90",x"FE",x"78", -- 0x3050
		x"6D",x"95",x"97",x"5A",x"D2",x"F0",x"E5",x"0F", -- 0x3058
		x"FF",x"DF",x"FF",x"DF",x"00",x"57",x"0F",x"DF", -- 0x3060
		x"E1",x"78",x"FF",x"55",x"04",x"55",x"F7",x"DD", -- 0x3068
		x"77",x"DD",x"77",x"FF",x"C3",x"FF",x"77",x"FF", -- 0x3070
		x"00",x"00",x"3C",x"87",x"78",x"F0",x"1E",x"F3", -- 0x3078
		x"B5",x"FF",x"D2",x"00",x"30",x"08",x"40",x"C2", -- 0x3080
		x"B0",x"4C",x"96",x"4A",x"95",x"D3",x"E7",x"DB", -- 0x3088
		x"EF",x"59",x"EF",x"4B",x"EF",x"F0",x"EF",x"33", -- 0x3090
		x"EF",x"48",x"EF",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x3098
		x"EF",x"3F",x"03",x"08",x"00",x"00",x"77",x"FF", -- 0x30A0
		x"77",x"FF",x"77",x"FF",x"77",x"DF",x"77",x"DF", -- 0x30A8
		x"00",x"57",x"0F",x"DF",x"F0",x"78",x"FF",x"55", -- 0x30B0
		x"00",x"55",x"FF",x"DD",x"FF",x"DD",x"FF",x"FF", -- 0x30B8
		x"67",x"7B",x"EF",x"7B",x"EF",x"6A",x"EF",x"7B", -- 0x30C0
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x30C8
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"CD",x"7B", -- 0x30D0
		x"FF",x"7B",x"EE",x"9D",x"FF",x"77",x"FF",x"FF", -- 0x30D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30F8
		x"FF",x"33",x"EE",x"1D",x"FF",x"7B",x"CD",x"7B", -- 0x3100
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3108
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3110
		x"EF",x"6A",x"EF",x"5B",x"67",x"5B",x"EF",x"5B", -- 0x3118
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3120
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3128
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3130
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3138
		x"EF",x"DB",x"EF",x"97",x"EF",x"D5",x"55",x"F3", -- 0x3140
		x"83",x"41",x"42",x"00",x"04",x"EE",x"19",x"FF", -- 0x3148
		x"19",x"FF",x"84",x"EE",x"84",x"00",x"C2",x"40", -- 0x3150
		x"C4",x"30",x"37",x"89",x"0C",x"01",x"0D",x"08", -- 0x3158
		x"FF",x"DD",x"FF",x"DD",x"00",x"55",x"4B",x"DD", -- 0x3160
		x"E1",x"78",x"F7",x"57",x"04",x"57",x"37",x"DF", -- 0x3168
		x"33",x"DF",x"71",x"FF",x"30",x"F7",x"97",x"FF", -- 0x3170
		x"E0",x"00",x"7C",x"87",x"B4",x"F0",x"DA",x"F3", -- 0x3178
		x"30",x"91",x"08",x"80",x"D1",x"40",x"00",x"02", -- 0x3180
		x"98",x"70",x"CC",x"B6",x"88",x"13",x"20",x"F3", -- 0x3188
		x"52",x"59",x"2B",x"4B",x"AB",x"F0",x"EB",x"33", -- 0x3190
		x"EF",x"48",x"EF",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x3198
		x"EF",x"3F",x"03",x"08",x"00",x"00",x"77",x"FF", -- 0x31A0
		x"55",x"FF",x"66",x"FF",x"77",x"DD",x"77",x"DD", -- 0x31A8
		x"00",x"55",x"0F",x"DD",x"F0",x"78",x"FF",x"57", -- 0x31B0
		x"00",x"57",x"FF",x"DF",x"FF",x"DF",x"FF",x"FF", -- 0x31B8
		x"67",x"7B",x"EF",x"7B",x"EF",x"6A",x"EF",x"7B", -- 0x31C0
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x31C8
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"CD",x"7B", -- 0x31D0
		x"FF",x"7B",x"EE",x"9D",x"FF",x"77",x"FF",x"FF", -- 0x31D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31F8
		x"FF",x"33",x"EE",x"1D",x"FF",x"7B",x"CD",x"7B", -- 0x3200
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3208
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3210
		x"EF",x"6A",x"EF",x"5B",x"67",x"5B",x"EF",x"5B", -- 0x3218
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3220
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3228
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3230
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3238
		x"EF",x"DB",x"EF",x"17",x"FE",x"00",x"40",x"40", -- 0x3240
		x"91",x"FF",x"77",x"FF",x"67",x"1F",x"CF",x"0F", -- 0x3248
		x"CF",x"0F",x"CF",x"0F",x"CF",x"0F",x"67",x"0F", -- 0x3250
		x"77",x"0F",x"33",x"1F",x"BB",x"FF",x"CC",x"FF", -- 0x3258
		x"FF",x"DF",x"FF",x"DF",x"00",x"57",x"83",x"DF", -- 0x3260
		x"01",x"78",x"B9",x"55",x"CC",x"55",x"FE",x"DD", -- 0x3268
		x"6E",x"D5",x"6E",x"77",x"6E",x"F7",x"4C",x"FF", -- 0x3270
		x"CC",x"00",x"DC",x"87",x"98",x"F0",x"12",x"F3", -- 0x3278
		x"80",x"C0",x"10",x"F0",x"88",x"40",x"4C",x"30", -- 0x3280
		x"AE",x"30",x"9F",x"30",x"FF",x"00",x"5D",x"33", -- 0x3288
		x"6E",x"71",x"DC",x"27",x"91",x"78",x"23",x"33", -- 0x3290
		x"EF",x"48",x"EF",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x3298
		x"67",x"3F",x"03",x"08",x"00",x"00",x"77",x"FF", -- 0x32A0
		x"77",x"77",x"77",x"FF",x"77",x"DB",x"77",x"DF", -- 0x32A8
		x"00",x"57",x"0F",x"DF",x"F0",x"78",x"FF",x"55", -- 0x32B0
		x"00",x"55",x"FF",x"DD",x"FF",x"DD",x"FF",x"FF", -- 0x32B8
		x"67",x"7B",x"EF",x"7B",x"EF",x"6A",x"EF",x"7B", -- 0x32C0
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x32C8
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"CD",x"7B", -- 0x32D0
		x"FF",x"7B",x"EE",x"9D",x"FF",x"77",x"FF",x"FF", -- 0x32D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x32F8
		x"FF",x"33",x"EE",x"1D",x"FF",x"7B",x"CD",x"7B", -- 0x3300
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3308
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3310
		x"EF",x"6A",x"EF",x"5B",x"67",x"5B",x"EF",x"5B", -- 0x3318
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3320
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3328
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3330
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3338
		x"EF",x"DB",x"DC",x"FE",x"99",x"FF",x"54",x"C0", -- 0x3340
		x"B0",x"30",x"D1",x"6E",x"22",x"3B",x"DD",x"B3", -- 0x3348
		x"44",x"51",x"80",x"60",x"AA",x"A0",x"DD",x"11", -- 0x3350
		x"F7",x"BF",x"E1",x"1E",x"B8",x"F0",x"A8",x"C0", -- 0x3358
		x"FF",x"DD",x"FF",x"DD",x"C8",x"55",x"CD",x"DD", -- 0x3360
		x"33",x"78",x"D1",x"DF",x"60",x"D7",x"EC",x"D7", -- 0x3368
		x"FC",x"D7",x"76",x"FF",x"75",x"FF",x"59",x"FF", -- 0x3370
		x"C0",x"00",x"B0",x"87",x"30",x"F0",x"9A",x"F3", -- 0x3378
		x"62",x"77",x"51",x"CC",x"00",x"00",x"40",x"00", -- 0x3380
		x"A9",x"4A",x"63",x"82",x"33",x"91",x"F7",x"33", -- 0x3388
		x"54",x"77",x"E8",x"CF",x"91",x"B8",x"22",x"33", -- 0x3390
		x"23",x"48",x"EF",x"5B",x"EF",x"5B",x"EF",x"5B", -- 0x3398
		x"67",x"3F",x"03",x"08",x"00",x"00",x"77",x"FF", -- 0x33A0
		x"77",x"77",x"77",x"FF",x"77",x"D9",x"77",x"DD", -- 0x33A8
		x"00",x"55",x"0F",x"DD",x"F0",x"78",x"FF",x"57", -- 0x33B0
		x"00",x"57",x"FF",x"DF",x"FF",x"DF",x"FF",x"FF", -- 0x33B8
		x"67",x"7B",x"EF",x"7B",x"EF",x"6A",x"EF",x"7B", -- 0x33C0
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x33C8
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"CD",x"7B", -- 0x33D0
		x"FF",x"7B",x"EE",x"9D",x"FF",x"77",x"FF",x"FF", -- 0x33D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33F8
		x"FF",x"33",x"EE",x"1D",x"FF",x"7B",x"CD",x"7B", -- 0x3400
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3408
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3410
		x"EF",x"6A",x"EF",x"5B",x"67",x"5B",x"EF",x"5B", -- 0x3418
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3420
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3428
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3430
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3438
		x"EF",x"60",x"FE",x"96",x"25",x"5B",x"99",x"CB", -- 0x3440
		x"01",x"3C",x"15",x"9D",x"47",x"4C",x"EF",x"A6", -- 0x3448
		x"EF",x"53",x"CF",x"D3",x"ED",x"1F",x"DC",x"5B", -- 0x3450
		x"3A",x"4B",x"0E",x"0F",x"F0",x"38",x"0F",x"0F", -- 0x3458
		x"FF",x"DF",x"33",x"DF",x"48",x"57",x"2D",x"DF", -- 0x3460
		x"E1",x"78",x"FF",x"55",x"00",x"55",x"77",x"DD", -- 0x3468
		x"77",x"DD",x"67",x"FF",x"67",x"F7",x"76",x"77", -- 0x3470
		x"02",x"00",x"0C",x"87",x"F0",x"F0",x"1E",x"F3", -- 0x3478
		x"BD",x"FE",x"03",x"68",x"00",x"A0",x"80",x"00", -- 0x3480
		x"40",x"4A",x"F7",x"53",x"FF",x"5B",x"EF",x"B9", -- 0x3488
		x"CD",x"59",x"CF",x"C9",x"BA",x"A2",x"24",x"45", -- 0x3490
		x"11",x"48",x"EF",x"4A",x"EF",x"5B",x"EF",x"5B", -- 0x3498
		x"E7",x"3F",x"01",x"08",x"00",x"00",x"77",x"FF", -- 0x34A0
		x"77",x"77",x"77",x"FF",x"77",x"DB",x"77",x"DF", -- 0x34A8
		x"00",x"57",x"0F",x"DF",x"F0",x"78",x"FF",x"55", -- 0x34B0
		x"08",x"55",x"FF",x"DD",x"FF",x"DD",x"FF",x"FF", -- 0x34B8
		x"67",x"7B",x"EF",x"7B",x"EF",x"6A",x"EF",x"7B", -- 0x34C0
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x34C8
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"CD",x"7B", -- 0x34D0
		x"FF",x"7B",x"EE",x"9D",x"FF",x"77",x"FF",x"FF", -- 0x34D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34F8
		x"FF",x"33",x"EE",x"1D",x"FF",x"7B",x"CD",x"7B", -- 0x3500
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3508
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x3510
		x"EF",x"6A",x"EF",x"5B",x"67",x"5B",x"EF",x"5B", -- 0x3518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3520
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3528
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3530
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3538
		x"EF",x"5B",x"EF",x"5B",x"23",x"5B",x"AB",x"4B", -- 0x3540
		x"44",x"F0",x"EF",x"33",x"EF",x"48",x"EF",x"4A", -- 0x3548
		x"EF",x"5B",x"AB",x"5B",x"67",x"5B",x"EF",x"5B", -- 0x3550
		x"23",x"4A",x"0C",x"0F",x"F0",x"30",x"0F",x"0D", -- 0x3558
		x"FF",x"DD",x"FF",x"DD",x"00",x"55",x"2D",x"DD", -- 0x3560
		x"E1",x"78",x"FF",x"57",x"00",x"57",x"77",x"DF", -- 0x3568
		x"77",x"DF",x"77",x"FF",x"77",x"FF",x"77",x"FF", -- 0x3570
		x"00",x"00",x"0C",x"87",x"F0",x"F0",x"96",x"F3", -- 0x3578
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3580
		x"CC",x"4A",x"FF",x"53",x"33",x"53",x"EE",x"1B", -- 0x3588
		x"CD",x"1B",x"CD",x"49",x"AB",x"68",x"67",x"48", -- 0x3590
		x"FF",x"48",x"EF",x"4A",x"EF",x"5B",x"EF",x"5B", -- 0x3598
		x"EF",x"3F",x"01",x"08",x"00",x"00",x"77",x"FF", -- 0x35A0
		x"77",x"FF",x"77",x"FF",x"77",x"DD",x"77",x"DD", -- 0x35A8
		x"00",x"55",x"0F",x"DD",x"F0",x"78",x"FF",x"57", -- 0x35B0
		x"08",x"57",x"FF",x"DF",x"FF",x"DF",x"FF",x"FF", -- 0x35B8
		x"67",x"7B",x"EF",x"7B",x"EF",x"6A",x"EF",x"7B", -- 0x35C0
		x"EF",x"7B",x"AB",x"7B",x"EF",x"7B",x"EF",x"7B", -- 0x35C8
		x"EF",x"7B",x"EF",x"7B",x"EF",x"7B",x"CD",x"7B", -- 0x35D0
		x"FF",x"7B",x"EE",x"9D",x"FF",x"77",x"FF",x"FF", -- 0x35D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3600
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3608
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3610
		x"FF",x"BC",x"FF",x"77",x"F0",x"E0",x"FF",x"FD", -- 0x3618
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x3620
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD", -- 0x3628
		x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"FF",x"77", -- 0x3630
		x"FF",x"66",x"FF",x"1F",x"F0",x"E1",x"FF",x"E7", -- 0x3638
		x"EF",x"ED",x"FF",x"00",x"FF",x"8B",x"FF",x"FF", -- 0x3640
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3658
		x"EE",x"4B",x"00",x"96",x"66",x"34",x"9E",x"D0", -- 0x3660
		x"FF",x"AC",x"FF",x"92",x"FE",x"ED",x"DF",x"CC", -- 0x3668
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x3670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3680
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3688
		x"FF",x"EF",x"FF",x"FE",x"FF",x"CE",x"FF",x"C8", -- 0x3690
		x"FF",x"08",x"FF",x"91",x"6C",x"73",x"CC",x"19", -- 0x3698
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"FF",x"FE", -- 0x36A0
		x"FF",x"FF",x"FE",x"77",x"EE",x"FF",x"FF",x"FF", -- 0x36A8
		x"FF",x"DC",x"EE",x"C8",x"7F",x"9A",x"13",x"10", -- 0x36B0
		x"20",x"DC",x"00",x"66",x"A8",x"D3",x"20",x"E7", -- 0x36B8
		x"FF",x"D0",x"FF",x"04",x"FF",x"9A",x"FF",x"FE", -- 0x36C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36D8
		x"42",x"0E",x"80",x"B4",x"E6",x"48",x"F8",x"80", -- 0x36E0
		x"DD",x"3B",x"FF",x"D1",x"FE",x"8C",x"FF",x"AC", -- 0x36E8
		x"BB",x"FA",x"DD",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x36F0
		x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x36F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3700
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x3708
		x"FF",x"88",x"FF",x"11",x"AA",x"77",x"EE",x"67", -- 0x3710
		x"EC",x"CF",x"C8",x"8F",x"E0",x"CF",x"EC",x"67", -- 0x3718
		x"FF",x"FF",x"FF",x"BB",x"FF",x"FF",x"DD",x"FF", -- 0x3720
		x"FF",x"FF",x"FF",x"EE",x"77",x"FC",x"33",x"EC", -- 0x3728
		x"21",x"E8",x"CC",x"D8",x"6E",x"50",x"3F",x"00", -- 0x3730
		x"3F",x"00",x"1F",x"31",x"3F",x"20",x"3F",x"20", -- 0x3738
		x"EE",x"33",x"FF",x"11",x"BB",x"A8",x"DD",x"EE", -- 0x3740
		x"FF",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3748
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3750
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3758
		x"6E",x"50",x"CC",x"00",x"30",x"33",x"C0",x"55", -- 0x3760
		x"CC",x"AE",x"EC",x"9F",x"EE",x"8F",x"FE",x"47", -- 0x3768
		x"FF",x"23",x"77",x"99",x"FF",x"FE",x"FF",x"FF", -- 0x3770
		x"FF",x"FF",x"EE",x"BB",x"FF",x"FF",x"FF",x"FF", -- 0x3778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EC",x"BB",x"80", -- 0x3788
		x"EE",x"11",x"EE",x"77",x"EC",x"FF",x"CC",x"FF", -- 0x3790
		x"D9",x"FF",x"C8",x"FF",x"40",x"77",x"C8",x"80", -- 0x3798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x37A0
		x"FF",x"FF",x"FF",x"EE",x"F3",x"FE",x"11",x"EC", -- 0x37A8
		x"CC",x"EC",x"EE",x"80",x"EE",x"51",x"CC",x"40", -- 0x37B0
		x"DC",x"00",x"DC",x"20",x"10",x"51",x"20",x"51", -- 0x37B8
		x"E8",x"60",x"EC",x"B8",x"FC",x"44",x"EE",x"77", -- 0x37C0
		x"FF",x"D1",x"77",x"EC",x"FF",x"FF",x"EC",x"FF", -- 0x37C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37D8
		x"40",x"D0",x"91",x"80",x"33",x"11",x"EE",x"00", -- 0x37E0
		x"99",x"A0",x"62",x"90",x"FE",x"70",x"EE",x"98", -- 0x37E8
		x"FF",x"EE",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF", -- 0x37F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3800
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"77", -- 0x3808
		x"EE",x"F3",x"DC",x"FE",x"FD",x"EE",x"FF",x"EC", -- 0x3810
		x"FD",x"DE",x"DB",x"45",x"38",x"78",x"11",x"73", -- 0x3818
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x3820
		x"FF",x"FF",x"FF",x"EE",x"D1",x"EF",x"BC",x"55", -- 0x3828
		x"EF",x"B3",x"7F",x"B3",x"B7",x"59",x"F7",x"63", -- 0x3830
		x"66",x"FB",x"CF",x"0F",x"86",x"38",x"34",x"0F", -- 0x3838
		x"DC",x"CD",x"FD",x"10",x"FF",x"8B",x"FF",x"3F", -- 0x3840
		x"FF",x"9E",x"FF",x"FC",x"FF",x"EE",x"FF",x"FF", -- 0x3848
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3850
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3858
		x"C0",x"3F",x"90",x"48",x"67",x"80",x"DE",x"00", -- 0x3860
		x"F0",x"10",x"C0",x"98",x"33",x"D5",x"FF",x"D5", -- 0x3868
		x"FF",x"73",x"FF",x"F9",x"FF",x"FF",x"FF",x"EE", -- 0x3870
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3878
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3880
		x"FF",x"FF",x"FF",x"FF",x"FC",x"7F",x"DB",x"FF", -- 0x3888
		x"BF",x"FE",x"FF",x"ED",x"FF",x"FF",x"FF",x"FF", -- 0x3890
		x"FF",x"88",x"FB",x"33",x"F0",x"85",x"DB",x"C4", -- 0x3898
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x38A0
		x"FF",x"FF",x"FF",x"EE",x"FF",x"FF",x"FF",x"DD", -- 0x38A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"FF",x"44", -- 0x38B0
		x"EE",x"FF",x"FF",x"0F",x"F0",x"F0",x"EF",x"C3", -- 0x38B8
		x"FD",x"E6",x"FD",x"00",x"FF",x"89",x"FF",x"FF", -- 0x38C0
		x"FF",x"FF",x"FF",x"DF",x"FF",x"FE",x"FF",x"FF", -- 0x38C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38D8
		x"75",x"3F",x"40",x"06",x"E2",x"00",x"FF",x"08", -- 0x38E0
		x"FF",x"08",x"EF",x"80",x"3C",x"DD",x"D1",x"DD", -- 0x38E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x38F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38F8
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"CF",x"F0", -- 0x3900
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3908
		x"CF",x"E0",x"CF",x"E0",x"CF",x"F0",x"CF",x"F0", -- 0x3910
		x"CF",x"F0",x"CF",x"F3",x"CF",x"F7",x"CF",x"F4", -- 0x3918
		x"FF",x"FF",x"FF",x"DF",x"FF",x"9D",x"F0",x"91", -- 0x3920
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"70",x"91", -- 0x3928
		x"B0",x"91",x"B0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3930
		x"F0",x"91",x"FE",x"91",x"FF",x"91",x"F1",x"91", -- 0x3938
		x"CF",x"F4",x"CF",x"F4",x"CF",x"F6",x"CF",x"F2", -- 0x3940
		x"CF",x"F0",x"CF",x"F7",x"CF",x"F7",x"CF",x"F1", -- 0x3948
		x"CF",x"F1",x"CF",x"F1",x"CF",x"F7",x"CF",x"F7", -- 0x3950
		x"CF",x"F0",x"CF",x"F7",x"CF",x"F7",x"CF",x"F0", -- 0x3958
		x"F1",x"91",x"F3",x"91",x"F2",x"91",x"F0",x"91", -- 0x3960
		x"F0",x"91",x"FC",x"91",x"FE",x"91",x"F3",x"91", -- 0x3968
		x"F1",x"91",x"F3",x"91",x"FE",x"91",x"FC",x"91", -- 0x3970
		x"F0",x"91",x"FF",x"91",x"FF",x"91",x"F9",x"91", -- 0x3978
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3980
		x"CF",x"F0",x"CF",x"F3",x"CF",x"F7",x"CF",x"F4", -- 0x3988
		x"CF",x"F4",x"CF",x"F4",x"CF",x"F6",x"CF",x"F2", -- 0x3990
		x"CF",x"F0",x"CF",x"F3",x"CF",x"F7",x"CF",x"F4", -- 0x3998
		x"F9",x"91",x"F9",x"91",x"FF",x"91",x"F6",x"91", -- 0x39A0
		x"F0",x"91",x"FE",x"91",x"FF",x"91",x"F1",x"91", -- 0x39A8
		x"F1",x"91",x"F3",x"91",x"F2",x"91",x"F0",x"91", -- 0x39B0
		x"F0",x"91",x"FE",x"91",x"FF",x"91",x"F1",x"91", -- 0x39B8
		x"CF",x"F4",x"CF",x"F4",x"CF",x"F7",x"CF",x"F3", -- 0x39C0
		x"CF",x"F0",x"CF",x"F7",x"CF",x"F7",x"CF",x"F0", -- 0x39C8
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F7",x"CF",x"F7", -- 0x39D0
		x"CF",x"F0",x"CF",x"0F",x"CF",x"0F",x"FF",x"FF", -- 0x39D8
		x"F1",x"91",x"F1",x"91",x"FF",x"91",x"FE",x"91", -- 0x39E0
		x"F0",x"91",x"FF",x"91",x"FF",x"91",x"F6",x"91", -- 0x39E8
		x"FC",x"91",x"F6",x"91",x"FF",x"91",x"FF",x"91", -- 0x39F0
		x"F0",x"91",x"0F",x"19",x"0F",x"1D",x"FF",x"FF", -- 0x39F8
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"CF",x"F0", -- 0x3A00
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3A08
		x"CF",x"E0",x"CF",x"E0",x"CF",x"F0",x"CF",x"F0", -- 0x3A10
		x"CF",x"F0",x"CF",x"F1",x"CF",x"F1",x"CF",x"F0", -- 0x3A18
		x"FF",x"FF",x"FF",x"DF",x"FF",x"9D",x"F0",x"91", -- 0x3A20
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"70",x"91", -- 0x3A28
		x"B0",x"91",x"B0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3A30
		x"F0",x"91",x"FC",x"91",x"FC",x"91",x"F0",x"91", -- 0x3A38
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3A40
		x"CF",x"F0",x"CF",x"F1",x"CF",x"F1",x"CF",x"F1", -- 0x3A48
		x"CF",x"F1",x"CF",x"F1",x"CF",x"F1",x"CF",x"F1", -- 0x3A50
		x"CF",x"F0",x"CF",x"F1",x"CF",x"F1",x"CF",x"F0", -- 0x3A58
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3A60
		x"F0",x"91",x"FC",x"91",x"FC",x"91",x"F0",x"91", -- 0x3A68
		x"F0",x"91",x"F0",x"91",x"FC",x"91",x"FC",x"91", -- 0x3A70
		x"F0",x"91",x"FC",x"91",x"FC",x"91",x"F8",x"91", -- 0x3A78
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3A80
		x"CF",x"F0",x"CF",x"F1",x"CF",x"F1",x"CF",x"F0", -- 0x3A88
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3A90
		x"CF",x"F0",x"CF",x"F1",x"CF",x"F1",x"CF",x"F0", -- 0x3A98
		x"F8",x"91",x"F8",x"91",x"FC",x"91",x"F4",x"91", -- 0x3AA0
		x"F0",x"91",x"FC",x"91",x"FC",x"91",x"F0",x"91", -- 0x3AA8
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3AB0
		x"F0",x"91",x"FC",x"91",x"FC",x"91",x"F0",x"91", -- 0x3AB8
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F1",x"CF",x"F1", -- 0x3AC0
		x"CF",x"F0",x"CF",x"F1",x"CF",x"F1",x"CF",x"F0", -- 0x3AC8
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F1",x"CF",x"F1", -- 0x3AD0
		x"CF",x"F0",x"CF",x"0F",x"CF",x"0F",x"FF",x"FF", -- 0x3AD8
		x"F0",x"91",x"F0",x"91",x"FC",x"91",x"FC",x"91", -- 0x3AE0
		x"F0",x"91",x"FC",x"91",x"FC",x"91",x"F4",x"91", -- 0x3AE8
		x"FC",x"91",x"F4",x"91",x"FC",x"91",x"FC",x"91", -- 0x3AF0
		x"F0",x"91",x"0F",x"19",x"0F",x"1D",x"FF",x"FF", -- 0x3AF8
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"CF",x"F0", -- 0x3B00
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B08
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B10
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B18
		x"FF",x"FF",x"FF",x"DF",x"FF",x"9D",x"F0",x"91", -- 0x3B20
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3B28
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3B30
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3B38
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B40
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B48
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B50
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B58
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3B60
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3B68
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3B70
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3B78
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B80
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B88
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B90
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3B98
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3BA0
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3BA8
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3BB0
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3BB8
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3BC0
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3BC8
		x"CF",x"F0",x"CF",x"F0",x"CF",x"F0",x"CF",x"F0", -- 0x3BD0
		x"CF",x"F0",x"CF",x"0F",x"CF",x"0F",x"FF",x"FF", -- 0x3BD8
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3BE0
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3BE8
		x"F0",x"91",x"F0",x"91",x"F0",x"91",x"F0",x"91", -- 0x3BF0
		x"F0",x"91",x"0F",x"19",x"0F",x"1D",x"FF",x"FF", -- 0x3BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C38
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3C40
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3C48
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3C50
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3C58
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3C60
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3C68
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3C70
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3C78
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3C80
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3C88
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3C90
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3C98
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3CA0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3CA8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3CB0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3CB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D38
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3D40
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3D48
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3D50
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3D58
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3D60
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3D68
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3D70
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3D78
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3D80
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3D88
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3D90
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3D98
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3DA0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3DA8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3DB0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3DB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E38
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3E40
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3E48
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3E50
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3E58
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3E60
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3E68
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3E70
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3E78
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3E80
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3E88
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3E90
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3E98
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3EA0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3EA8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3EB0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3ED8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F38
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3F40
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3F48
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3F50
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3F58
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3F60
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3F68
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3F70
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x3F78
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3F80
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3F88
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3F90
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3F98
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3FA0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3FA8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3FB0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x3FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
