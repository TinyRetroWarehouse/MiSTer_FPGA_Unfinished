-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_A5 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_A5 is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"FB",x"FF",x"EF",x"C3",x"61",x"31",x"9B",x"1A", -- 0x0000
		x"5E",x"7F",x"8F",x"47",x"03",x"20",x"31",x"11", -- 0x0008
		x"FF",x"FB",x"FF",x"FF",x"F7",x"F3",x"31",x"99", -- 0x0010
		x"1D",x"9F",x"FF",x"FF",x"1F",x"23",x"31",x"98", -- 0x0018
		x"7E",x"3F",x"BF",x"3F",x"47",x"22",x"24",x"46", -- 0x0020
		x"03",x"40",x"A8",x"A9",x"8C",x"66",x"54",x"B0", -- 0x0028
		x"FF",x"FF",x"FF",x"F7",x"FF",x"7F",x"3D",x"3F", -- 0x0030
		x"1E",x"B8",x"73",x"0D",x"A2",x"30",x"56",x"0C", -- 0x0038
		x"FF",x"3F",x"9B",x"01",x"09",x"5B",x"4C",x"38", -- 0x0040
		x"28",x"2C",x"04",x"B7",x"05",x"15",x"88",x"40", -- 0x0048
		x"FF",x"3F",x"1F",x"BF",x"FF",x"FF",x"FF",x"7F", -- 0x0050
		x"7F",x"CF",x"87",x"47",x"67",x"3B",x"97",x"30", -- 0x0058
		x"7F",x"FF",x"9F",x"9F",x"0E",x"9C",x"BC",x"42", -- 0x0060
		x"22",x"41",x"91",x"CB",x"6E",x"20",x"00",x"10", -- 0x0068
		x"FF",x"FF",x"FF",x"EF",x"C7",x"D7",x"67",x"3F", -- 0x0070
		x"7D",x"FF",x"FF",x"CF",x"C7",x"67",x"3F",x"7F", -- 0x0078
		x"FF",x"BF",x"FF",x"E7",x"53",x"23",x"23",x"BF", -- 0x0080
		x"7F",x"7E",x"90",x"A0",x"90",x"69",x"50",x"B0", -- 0x0088
		x"FF",x"FF",x"EF",x"FF",x"FF",x"FB",x"F9",x"F9", -- 0x0090
		x"CF",x"87",x"E3",x"43",x"67",x"E7",x"FF",x"FF", -- 0x0098
		x"20",x"48",x"C5",x"83",x"45",x"A8",x"08",x"09", -- 0x00A0
		x"05",x"68",x"B4",x"0D",x"06",x"02",x"21",x"11", -- 0x00A8
		x"FF",x"F3",x"E1",x"D9",x"51",x"08",x"AD",x"73", -- 0x00B0
		x"7B",x"FB",x"BF",x"1F",x"BF",x"2B",x"11",x"19", -- 0x00B8
		x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"F1",x"F3", -- 0x00C0
		x"F9",x"FF",x"FF",x"FB",x"D0",x"D8",x"A1",x"11", -- 0x00C8
		x"FF",x"FF",x"FF",x"FF",x"BF",x"1F",x"1F",x"BF", -- 0x00D0
		x"DE",x"F4",x"F8",x"EC",x"1D",x"2A",x"20",x"18", -- 0x00D8
		x"FF",x"BF",x"FF",x"FF",x"F8",x"E8",x"E8",x"B0", -- 0x00E0
		x"04",x"14",x"0A",x"B3",x"09",x"15",x"8B",x"41", -- 0x00E8
		x"FC",x"F0",x"E8",x"C6",x"E1",x"80",x"10",x"40", -- 0x00F0
		x"35",x"A2",x"C8",x"B0",x"A4",x"B9",x"D6",x"30", -- 0x00F8
		x"EF",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0100
		x"FC",x"FB",x"EA",x"F1",x"E5",x"D1",x"40",x"F0", -- 0x0108
		x"FE",x"FE",x"FC",x"F2",x"E1",x"B8",x"90",x"5A", -- 0x0110
		x"4B",x"20",x"74",x"E0",x"70",x"89",x"56",x"30", -- 0x0118
		x"FF",x"FE",x"FE",x"EC",x"C3",x"C7",x"EF",x"E7", -- 0x0120
		x"F3",x"FF",x"FF",x"FF",x"FF",x"FE",x"FD",x"F9", -- 0x0128
		x"FC",x"78",x"32",x"32",x"51",x"D8",x"CA",x"D1", -- 0x0130
		x"A5",x"C6",x"6B",x"75",x"D2",x"88",x"86",x"44", -- 0x0138
		x"FF",x"DF",x"FF",x"FF",x"F7",x"C2",x"A2",x"B1", -- 0x0140
		x"21",x"33",x"1F",x"0F",x"9F",x"FF",x"FF",x"FC", -- 0x0148
		x"FF",x"F9",x"FC",x"EF",x"57",x"67",x"3F",x"7F", -- 0x0150
		x"FD",x"FE",x"F7",x"F5",x"E2",x"A0",x"76",x"E4", -- 0x0158
		x"FF",x"CE",x"FE",x"FE",x"FF",x"FF",x"FA",x"E8", -- 0x0160
		x"F1",x"D8",x"D4",x"FD",x"8F",x"92",x"81",x"D1", -- 0x0168
		x"A0",x"98",x"D4",x"40",x"20",x"42",x"28",x"94", -- 0x0170
		x"58",x"58",x"08",x"A4",x"95",x"2A",x"20",x"18", -- 0x0178
		x"60",x"08",x"AA",x"50",x"78",x"14",x"8B",x"CF", -- 0x0180
		x"3F",x"FC",x"FC",x"F4",x"F2",x"FB",x"F9",x"FF", -- 0x0188
		x"31",x"4D",x"A3",x"3F",x"BF",x"FF",x"E7",x"E3", -- 0x0190
		x"A3",x"97",x"DF",x"7F",x"7F",x"7F",x"FF",x"FF", -- 0x0198
		x"E0",x"30",x"93",x"04",x"05",x"56",x"42",x"23", -- 0x01A0
		x"21",x"0E",x"06",x"AF",x"1F",x"9F",x"FF",x"FF", -- 0x01A8
		x"10",x"44",x"24",x"96",x"93",x"DA",x"52",x"41", -- 0x01B0
		x"77",x"A3",x"63",x"77",x"3F",x"0F",x"FF",x"FF", -- 0x01B8
		x"D1",x"B8",x"E8",x"E1",x"22",x"86",x"82",x"C3", -- 0x01C0
		x"69",x"04",x"97",x"CE",x"8C",x"9C",x"FE",x"FF", -- 0x01C8
		x"A6",x"41",x"41",x"2B",x"3B",x"1F",x"9F",x"1F", -- 0x01D0
		x"BF",x"67",x"E3",x"E3",x"23",x"73",x"77",x"7F", -- 0x01D8
		x"10",x"B8",x"ED",x"EF",x"37",x"8E",x"82",x"47", -- 0x01E0
		x"6F",x"27",x"8F",x"CF",x"8E",x"DC",x"7C",x"3E", -- 0x01E8
		x"FF",x"FF",x"EF",x"F7",x"67",x"23",x"77",x"3F", -- 0x01F0
		x"FF",x"FF",x"CF",x"87",x"C7",x"67",x"7F",x"7F", -- 0x01F8
		x"11",x"B9",x"E9",x"AF",x"17",x"87",x"CF",x"FE", -- 0x0200
		x"32",x"71",x"F9",x"CF",x"C7",x"EF",x"FC",x"FC", -- 0x0208
		x"FF",x"FF",x"CF",x"87",x"C7",x"A7",x"FF",x"7F", -- 0x0210
		x"1F",x"3F",x"FD",x"FC",x"3F",x"9F",x"FF",x"7F", -- 0x0218
		x"E0",x"28",x"8D",x"05",x"07",x"43",x"4F",x"2E", -- 0x0220
		x"24",x"0C",x"08",x"A2",x"08",x"05",x"85",x"41", -- 0x0228
		x"0B",x"6F",x"A7",x"67",x"47",x"67",x"BF",x"6F", -- 0x0230
		x"2F",x"BF",x"1F",x"3F",x"3F",x"3D",x"7D",x"FF", -- 0x0238
		x"C0",x"20",x"92",x"9C",x"C9",x"DF",x"EE",x"FF", -- 0x0240
		x"FF",x"FD",x"F8",x"E8",x"C5",x"CF",x"FF",x"FF", -- 0x0248
		x"08",x"54",x"24",x"1A",x"AD",x"FA",x"D0",x"39", -- 0x0250
		x"DC",x"C3",x"E7",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x0258
		x"11",x"B8",x"6A",x"EF",x"35",x"8E",x"84",x"C4", -- 0x0260
		x"6A",x"3F",x"F3",x"F9",x"FF",x"FF",x"FD",x"FC", -- 0x0268
		x"E6",x"41",x"00",x"20",x"E8",x"B9",x"13",x"0D", -- 0x0270
		x"A2",x"F9",x"B1",x"9C",x"0C",x"8A",x"27",x"F1", -- 0x0278
		x"B0",x"49",x"A8",x"CF",x"F4",x"EE",x"D7",x"63", -- 0x0280
		x"25",x"91",x"D1",x"62",x"B3",x"2F",x"AF",x"FF", -- 0x0288
		x"A0",x"98",x"D4",x"C0",x"A0",x"42",x"08",x"84", -- 0x0290
		x"00",x"A0",x"D0",x"EC",x"8D",x"D6",x"FB",x"FD", -- 0x0298
		x"FF",x"FE",x"FF",x"FE",x"FE",x"FC",x"FE",x"F7", -- 0x02A0
		x"F4",x"F4",x"F2",x"F9",x"FD",x"FD",x"FD",x"FF", -- 0x02A8
		x"68",x"74",x"24",x"5A",x"DD",x"36",x"48",x"2C", -- 0x02B0
		x"2D",x"FA",x"3E",x"32",x"7B",x"FB",x"FD",x"FD", -- 0x02B8
		x"FE",x"9E",x"9F",x"FF",x"FB",x"F9",x"E9",x"EF", -- 0x02C0
		x"E7",x"FF",x"FE",x"FA",x"FF",x"D3",x"F9",x"FF", -- 0x02C8
		x"B6",x"CC",x"7A",x"DE",x"DD",x"EC",x"F6",x"9F", -- 0x02D0
		x"0D",x"47",x"23",x"73",x"1F",x"BF",x"FF",x"FF", -- 0x02D8
		x"A0",x"41",x"4B",x"BD",x"F3",x"B0",x"D8",x"E8", -- 0x02E0
		x"F0",x"DA",x"CC",x"FD",x"CF",x"F2",x"F8",x"FE", -- 0x02E8
		x"A0",x"98",x"D4",x"C0",x"A0",x"EA",x"34",x"90", -- 0x02F0
		x"60",x"48",x"48",x"C4",x"C5",x"A2",x"A0",x"D8", -- 0x02F8
		x"FE",x"DF",x"CA",x"FF",x"F4",x"F3",x"FB",x"F8", -- 0x0300
		x"FF",x"FE",x"FE",x"FF",x"FD",x"FD",x"FC",x"FA", -- 0x0308
		x"A0",x"18",x"14",x"20",x"10",x"1A",x"C8",x"F4", -- 0x0310
		x"60",x"88",x"88",x"64",x"95",x"8A",x"A0",x"D8", -- 0x0318
		x"20",x"40",x"CA",x"89",x"47",x"A8",x"12",x"09", -- 0x0320
		x"29",x"4C",x"AC",x"15",x"06",x"12",x"21",x"11", -- 0x0328
		x"FF",x"7F",x"FF",x"FF",x"BF",x"1E",x"9D",x"3F", -- 0x0330
		x"BF",x"BF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF", -- 0x0338
		x"11",x"B0",x"EC",x"EB",x"32",x"88",x"CE",x"F9", -- 0x0340
		x"74",x"B3",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0348
		x"E6",x"C1",x"C0",x"20",x"28",x"15",x"1F",x"0D", -- 0x0350
		x"6E",x"FF",x"FF",x"BF",x"3F",x"FF",x"FF",x"FF", -- 0x0358
		x"DF",x"CF",x"FF",x"FF",x"FF",x"F7",x"F3",x"D9", -- 0x0360
		x"50",x"28",x"0A",x"13",x"9C",x"8C",x"45",x"12", -- 0x0368
		x"FF",x"FF",x"FF",x"FF",x"DF",x"CF",x"0F",x"85", -- 0x0370
		x"A4",x"C4",x"75",x"32",x"68",x"46",x"8B",x"80", -- 0x0378
		x"FF",x"FE",x"F2",x"E1",x"B3",x"23",x"34",x"18", -- 0x0380
		x"94",x"8E",x"C7",x"E3",x"D5",x"D9",x"97",x"CF", -- 0x0388
		x"FF",x"7F",x"FF",x"F9",x"FC",x"FF",x"FF",x"7F", -- 0x0390
		x"7F",x"FF",x"FF",x"D3",x"EB",x"B1",x"1B",x"8F", -- 0x0398
		x"FF",x"FF",x"FE",x"FC",x"F6",x"F3",x"F1",x"F1", -- 0x03A0
		x"F7",x"CE",x"CF",x"FF",x"FF",x"9F",x"FF",x"FF", -- 0x03A8
		x"FF",x"FB",x"6D",x"E1",x"34",x"88",x"10",x"3B", -- 0x03B0
		x"0F",x"8F",x"DF",x"F7",x"F3",x"CD",x"CF",x"FF", -- 0x03B8
		x"11",x"B8",x"E8",x"EE",x"34",x"8D",x"86",x"C4", -- 0x03C0
		x"6E",x"87",x"C3",x"C1",x"E3",x"FF",x"FF",x"FF", -- 0x03C8
		x"E6",x"C1",x"C0",x"20",x"A8",x"19",x"13",x"0D", -- 0x03D0
		x"A2",x"F9",x"B1",x"1C",x"0C",x"8A",x"C7",x"F9", -- 0x03D8
		x"C0",x"20",x"12",x"9C",x"09",x"1E",x"8C",x"CE", -- 0x03E0
		x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03E8
		x"08",x"54",x"64",x"5A",x"ED",x"FA",x"D0",x"39", -- 0x03F0
		x"1C",x"0F",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03F8
		x"11",x"B8",x"E8",x"EE",x"34",x"8D",x"C6",x"E0", -- 0x0400
		x"6C",x"07",x"83",x"C3",x"F7",x"FF",x"FF",x"FF", -- 0x0408
		x"E6",x"C1",x"C0",x"20",x"A8",x"15",x"1F",x"0D", -- 0x0410
		x"04",x"C6",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0418
		x"60",x"38",x"92",x"60",x"68",x"30",x"B8",x"C9", -- 0x0420
		x"1F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0428
		x"31",x"4D",x"C7",x"67",x"EF",x"FF",x"FF",x"FF", -- 0x0430
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0438
		x"20",x"41",x"C8",x"89",x"47",x"A8",x"10",x"09", -- 0x0440
		x"11",x"58",x"AC",x"5D",x"2E",x"12",x"21",x"11", -- 0x0448
		x"A0",x"98",x"D4",x"C0",x"A0",x"C2",x"28",x"14", -- 0x0450
		x"00",x"88",x"88",x"24",x"95",x"2A",x"20",x"18", -- 0x0458
		x"62",x"20",x"92",x"61",x"4A",x"20",x"26",x"51", -- 0x0460
		x"88",x"44",x"AE",x"AB",x"98",x"66",x"58",x"B0", -- 0x0468
		x"36",x"4C",x"D2",x"22",x"51",x"38",x"8A",x"B9", -- 0x0470
		x"D5",x"86",x"2B",x"B5",x"92",x"88",x"86",x"44", -- 0x0478
		x"C0",x"20",x"93",x"0C",x"05",x"52",x"44",x"28", -- 0x0480
		x"20",x"1A",x"0E",x"B3",x"0D",x"15",x"88",x"40", -- 0x0488
		x"08",x"54",x"24",x"9A",x"AD",x"FA",x"50",x"20", -- 0x0490
		x"15",x"A2",x"E0",x"D0",x"64",x"F9",x"56",x"30", -- 0x0498
		x"11",x"B8",x"E8",x"EE",x"34",x"8D",x"86",x"40", -- 0x04A0
		x"6C",x"07",x"92",x"C9",x"8D",x"C0",x"40",x"10", -- 0x04A8
		x"E6",x"C1",x"C0",x"20",x"A8",x"19",x"13",x"0D", -- 0x04B0
		x"82",x"29",x"19",x"04",x"18",x"86",x"CB",x"00", -- 0x04B8
		x"7B",x"D6",x"AD",x"FF",x"B7",x"DF",x"7E",x"DF", -- 0x04C0
		x"FF",x"FF",x"FB",x"FE",x"BF",x"FF",x"EF",x"7B", -- 0x04C8
		x"FF",x"FF",x"DF",x"DF",x"FD",x"FF",x"F7",x"FF", -- 0x04D0
		x"BB",x"FD",x"FF",x"FF",x"FF",x"FD",x"BF",x"EF", -- 0x04D8
		x"FF",x"FF",x"DB",x"F7",x"DF",x"FB",x"BF",x"FF", -- 0x04E0
		x"F9",x"ED",x"FE",x"DD",x"B3",x"FF",x"FD",x"DF", -- 0x04E8
		x"7F",x"DB",x"EF",x"FD",x"D9",x"CB",x"BF",x"5F", -- 0x04F0
		x"B3",x"FD",x"F2",x"F6",x"BD",x"FD",x"FF",x"FF", -- 0x04F8
		x"FF",x"FD",x"FF",x"FF",x"DF",x"FF",x"F7",x"FE", -- 0x0500
		x"FF",x"FE",x"FE",x"FF",x"FF",x"FD",x"FF",x"FF", -- 0x0508
		x"67",x"BB",x"F7",x"ED",x"7E",x"6B",x"BF",x"5F", -- 0x0510
		x"EB",x"7F",x"9F",x"DB",x"F9",x"FF",x"FF",x"FF", -- 0x0518
		x"9F",x"DE",x"E7",x"C3",x"DF",x"DC",x"8D",x"BB", -- 0x0520
		x"DB",x"EF",x"FF",x"FF",x"FF",x"E7",x"F3",x"FF", -- 0x0528
		x"FF",x"FD",x"FD",x"DF",x"6F",x"7F",x"23",x"EC", -- 0x0530
		x"E7",x"D7",x"D7",x"CF",x"ED",x"BD",x"9F",x"FF", -- 0x0538
		x"BF",x"9F",x"FF",x"FF",x"FB",x"E1",x"EF",x"CE", -- 0x0540
		x"FD",x"DE",x"EC",x"DF",x"FB",x"F5",x"FF",x"FF", -- 0x0548
		x"FF",x"FF",x"BF",x"DD",x"FD",x"FF",x"FF",x"DF", -- 0x0550
		x"7F",x"DF",x"EB",x"67",x"EF",x"7B",x"FE",x"EF", -- 0x0558
		x"FF",x"EF",x"DF",x"FF",x"FF",x"DB",x"97",x"2F", -- 0x0560
		x"B9",x"DE",x"9E",x"8F",x"FF",x"FB",x"F7",x"FF", -- 0x0568
		x"FF",x"FF",x"7D",x"AF",x"BF",x"FB",x"F7",x"7F", -- 0x0570
		x"E7",x"BB",x"3F",x"D7",x"EF",x"E3",x"DC",x"FF", -- 0x0578
		x"BF",x"DF",x"FE",x"FE",x"EE",x"BF",x"B3",x"F7", -- 0x0580
		x"D7",x"FD",x"79",x"9F",x"C7",x"DF",x"BB",x"FD", -- 0x0588
		x"DF",x"67",x"FF",x"BF",x"6F",x"7F",x"EF",x"FF", -- 0x0590
		x"BF",x"DF",x"FB",x"AB",x"BF",x"FF",x"FF",x"FF", -- 0x0598
		x"DF",x"FD",x"FE",x"F3",x"FB",x"E7",x"75",x"AF", -- 0x05A0
		x"CD",x"F6",x"C6",x"9D",x"FF",x"59",x"BD",x"FF", -- 0x05A8
		x"FE",x"FE",x"FF",x"BF",x"FF",x"FF",x"DF",x"B7", -- 0x05B0
		x"DF",x"CB",x"BF",x"EF",x"FF",x"7F",x"BB",x"1F", -- 0x05B8
		x"FF",x"FC",x"DB",x"F7",x"FD",x"F9",x"F7",x"FF", -- 0x05C0
		x"FD",x"FD",x"FE",x"DD",x"FB",x"ED",x"FF",x"FF", -- 0x05C8
		x"7F",x"DF",x"AF",x"1D",x"BD",x"CB",x"BF",x"DF", -- 0x05D0
		x"A3",x"2D",x"72",x"76",x"BD",x"FD",x"FC",x"FF", -- 0x05D8
		x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x05E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F8
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x0600
		x"FF",x"FF",x"FF",x"DF",x"FB",x"FF",x"FF",x"FF", -- 0x0608
		x"FF",x"EF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FB", -- 0x0610
		x"F7",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x0618
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"DF",x"FF", -- 0x0620
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0628
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0630
		x"FF",x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x0638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0640
		x"FF",x"FE",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF", -- 0x0648
		x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"FF",x"FF", -- 0x0650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0658
		x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x0660
		x"F9",x"64",x"98",x"98",x"8C",x"0F",x"0B",x"BF", -- 0x0668
		x"FF",x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF", -- 0x0670
		x"FF",x"FB",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF", -- 0x0678
		x"FF",x"EF",x"FF",x"DF",x"FF",x"FF",x"BF",x"FF", -- 0x0680
		x"FF",x"FF",x"FE",x"FE",x"BC",x"F8",x"FC",x"FE", -- 0x0688
		x"FF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0690
		x"BF",x"F9",x"F0",x"78",x"10",x"3A",x"7F",x"3F", -- 0x0698
		x"FB",x"FD",x"FC",x"DC",x"58",x"0E",x"9D",x"0E", -- 0x06A0
		x"0F",x"9F",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x06A8
		x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"FF",x"7D", -- 0x06B0
		x"FF",x"FF",x"FF",x"EF",x"F7",x"7F",x"FF",x"FF", -- 0x06B8
		x"FF",x"FB",x"FF",x"FD",x"F8",x"F8",x"D8",x"FC", -- 0x06C0
		x"FF",x"FF",x"FF",x"FB",x"DF",x"FF",x"FF",x"FD", -- 0x06C8
		x"FF",x"E7",x"E3",x"73",x"63",x"EB",x"77",x"FF", -- 0x06D0
		x"FF",x"BF",x"FF",x"FF",x"FF",x"FB",x"FF",x"FF", -- 0x06D8
		x"FF",x"FF",x"7D",x"6E",x"79",x"FF",x"4F",x"FE", -- 0x06E0
		x"FD",x"79",x"B6",x"FF",x"EF",x"6F",x"F7",x"FF", -- 0x06E8
		x"9F",x"B7",x"B5",x"FF",x"FB",x"FD",x"FF",x"7E", -- 0x06F0
		x"D7",x"FF",x"FF",x"CF",x"FE",x"BC",x"FB",x"E3", -- 0x06F8
		x"FD",x"F7",x"DB",x"DE",x"FD",x"FB",x"F7",x"BF", -- 0x0700
		x"B7",x"FB",x"F7",x"FF",x"FB",x"C9",x"B1",x"FB", -- 0x0708
		x"FF",x"FF",x"FF",x"77",x"BF",x"FF",x"BB",x"CE", -- 0x0710
		x"EF",x"69",x"D7",x"FD",x"AD",x"8F",x"FF",x"FF", -- 0x0718
		x"BE",x"BF",x"FE",x"ED",x"DF",x"FF",x"7F",x"FF", -- 0x0720
		x"FF",x"FF",x"B7",x"FF",x"FD",x"EF",x"FB",x"FB", -- 0x0728
		x"F7",x"FB",x"FB",x"8F",x"AF",x"79",x"3D",x"B6", -- 0x0730
		x"C4",x"FF",x"FF",x"FF",x"F9",x"BB",x"73",x"FF", -- 0x0738
		x"FF",x"FF",x"F7",x"FF",x"DB",x"FF",x"FF",x"FF", -- 0x0740
		x"FF",x"FF",x"FF",x"F7",x"DF",x"FF",x"FF",x"FF", -- 0x0748
		x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"7F",x"FB", -- 0x0750
		x"F7",x"FF",x"BF",x"EF",x"FF",x"FF",x"FB",x"FF", -- 0x0758
		x"DF",x"FF",x"F7",x"FF",x"DB",x"FF",x"FF",x"FF", -- 0x0760
		x"FF",x"FF",x"FF",x"F7",x"DF",x"FF",x"FF",x"FF", -- 0x0768
		x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"7F",x"FB", -- 0x0770
		x"F7",x"FF",x"BF",x"EF",x"FF",x"FF",x"FB",x"FF", -- 0x0778
		x"FF",x"FF",x"FF",x"DE",x"FF",x"FF",x"FF",x"FF", -- 0x0780
		x"EF",x"FF",x"FF",x"FF",x"FD",x"FF",x"DF",x"FF", -- 0x0788
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB", -- 0x0790
		x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x0798
		x"FF",x"FF",x"FF",x"FE",x"FF",x"DF",x"FF",x"FD", -- 0x07A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"FF", -- 0x07A8
		x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB", -- 0x07B0
		x"FF",x"FF",x"BD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B8
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"FF",x"EF", -- 0x07C0
		x"FF",x"FE",x"F7",x"F7",x"DF",x"FF",x"DF",x"FF", -- 0x07C8
		x"FF",x"7F",x"FF",x"EF",x"EF",x"FF",x"FF",x"FB", -- 0x07D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FF", -- 0x07D8
		x"FF",x"BF",x"FF",x"FF",x"FF",x"DF",x"FD",x"FF", -- 0x07E0
		x"FB",x"DF",x"DF",x"F7",x"FB",x"BF",x"FF",x"FF", -- 0x07E8
		x"FF",x"7F",x"EF",x"FF",x"AF",x"FF",x"FB",x"FB", -- 0x07F0
		x"FD",x"DF",x"FF",x"FF",x"F7",x"F7",x"FB",x"FF", -- 0x07F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0800
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0808
		x"F7",x"7B",x"BF",x"BF",x"BF",x"FF",x"DF",x"DD", -- 0x0810
		x"CF",x"EF",x"F7",x"F7",x"FB",x"FB",x"F9",x"FC", -- 0x0818
		x"7F",x"B7",x"BF",x"CF",x"FF",x"FF",x"F7",x"FB", -- 0x0820
		x"FB",x"FF",x"FD",x"FE",x"FE",x"FE",x"FF",x"FF", -- 0x0828
		x"FF",x"F7",x"FB",x"F7",x"FF",x"DF",x"FF",x"FF", -- 0x0830
		x"FF",x"EF",x"FF",x"FD",x"AD",x"FF",x"FF",x"7F", -- 0x0838
		x"FF",x"FE",x"FF",x"FE",x"FE",x"FF",x"FF",x"FF", -- 0x0840
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0848
		x"7F",x"FD",x"FB",x"FF",x"F7",x"7F",x"FF",x"3F", -- 0x0850
		x"3F",x"7F",x"F9",x"7D",x"3B",x"7F",x"FF",x"7F", -- 0x0858
		x"FF",x"ED",x"EF",x"FF",x"FF",x"FF",x"DF",x"3F", -- 0x0860
		x"9D",x"E4",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0868
		x"FF",x"FF",x"F7",x"FF",x"FF",x"BF",x"7F",x"BF", -- 0x0870
		x"F7",x"FB",x"EF",x"7F",x"BF",x"E7",x"F9",x"FE", -- 0x0878
		x"FF",x"FF",x"EC",x"FF",x"FF",x"FF",x"5E",x"7F", -- 0x0880
		x"DB",x"E7",x"FB",x"FD",x"FF",x"FE",x"FE",x"FF", -- 0x0888
		x"FF",x"77",x"77",x"FF",x"FF",x"FF",x"FF",x"FD", -- 0x0890
		x"FD",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x0898
		x"FF",x"DF",x"DF",x"FE",x"F7",x"BF",x"9E",x"49", -- 0x08A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08A8
		x"FF",x"FB",x"DF",x"DF",x"6F",x"7F",x"7F",x"7C", -- 0x08B0
		x"9B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08B8
		x"7F",x"9B",x"E3",x"FC",x"FE",x"FF",x"FF",x"FF", -- 0x08C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08C8
		x"FF",x"7D",x"FF",x"FF",x"7F",x"8F",x"F3",x"F9", -- 0x08D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08E8
		x"7F",x"2F",x"AB",x"CF",x"FF",x"FA",x"F9",x"FF", -- 0x08F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08F8
		x"76",x"AF",x"CB",x"F7",x"FB",x"FD",x"FC",x"FF", -- 0x0900
		x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0908
		x"FF",x"6F",x"EF",x"BB",x"F9",x"7F",x"FD",x"DF", -- 0x0910
		x"DF",x"0F",x"CF",x"EB",x"FB",x"FB",x"FD",x"FE", -- 0x0918
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0920
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0928
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0930
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0938
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0940
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0948
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0950
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0958
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0960
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0968
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0978
		x"7F",x"F7",x"BF",x"CF",x"DF",x"FF",x"DF",x"CB", -- 0x0980
		x"DF",x"CF",x"ED",x"E7",x"EB",x"F7",x"FF",x"F7", -- 0x0988
		x"FF",x"F7",x"FB",x"77",x"7F",x"BF",x"FF",x"FF", -- 0x0990
		x"FF",x"EF",x"FF",x"FD",x"AD",x"FF",x"FF",x"7F", -- 0x0998
		x"FF",x"F7",x"FF",x"F9",x"FB",x"FD",x"FD",x"FE", -- 0x09A0
		x"FD",x"FF",x"FF",x"FE",x"FE",x"FF",x"FF",x"FF", -- 0x09A8
		x"7F",x"FD",x"FB",x"FF",x"F7",x"7F",x"FF",x"FF", -- 0x09B0
		x"FF",x"7F",x"F9",x"7D",x"3B",x"7F",x"FF",x"7F", -- 0x09B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09C8
		x"F7",x"7B",x"3F",x"BF",x"BF",x"BF",x"DF",x"D9", -- 0x09D0
		x"ED",x"DF",x"FF",x"E7",x"EB",x"EF",x"F7",x"F6", -- 0x09D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09E8
		x"F7",x"FB",x"F3",x"FF",x"FB",x"FF",x"FD",x"F9", -- 0x09F0
		x"FF",x"FD",x"FF",x"FD",x"FC",x"FF",x"FF",x"FE", -- 0x09F8
		x"F6",x"FF",x"FB",x"FB",x"FD",x"FF",x"FE",x"FF", -- 0x0A00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A08
		x"FF",x"6F",x"EF",x"BB",x"F9",x"7F",x"FD",x"DF", -- 0x0A10
		x"DF",x"8F",x"CF",x"EB",x"FB",x"FB",x"FD",x"FE", -- 0x0A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A28
		x"FF",x"F5",x"EB",x"EF",x"F7",x"EF",x"FF",x"EF", -- 0x0A30
		x"F7",x"F7",x"F9",x"ED",x"FF",x"FF",x"EF",x"FF", -- 0x0A38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A58
		x"C7",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC", -- 0x0A60
		x"FC",x"FC",x"FC",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x0A68
		x"07",x"07",x"0F",x"0F",x"07",x"07",x"07",x"17", -- 0x0A70
		x"11",x"1F",x"0F",x"0F",x"07",x"3F",x"3F",x"3F", -- 0x0A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x0A80
		x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A88
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",x"00", -- 0x0A90
		x"00",x"00",x"00",x"F0",x"F0",x"F0",x"FE",x"FE", -- 0x0A98
		x"FF",x"FF",x"FF",x"3F",x"3F",x"3F",x"3F",x"3F", -- 0x0AA0
		x"3F",x"03",x"03",x"03",x"03",x"03",x"07",x"FF", -- 0x0AA8
		x"FE",x"F8",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x0AB0
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"FE", -- 0x0AB8
		x"FF",x"FF",x"FF",x"F0",x"E0",x"E0",x"E0",x"F1", -- 0x0AC0
		x"F1",x"F1",x"F1",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x0AC8
		x"FE",x"F8",x"F0",x"00",x"00",x"00",x"00",x"F0", -- 0x0AD0
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"FE", -- 0x0AD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"0E",x"0E", -- 0x0AE0
		x"0E",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x0AE8
		x"FE",x"E0",x"C0",x"C0",x"C0",x"00",x"00",x"00", -- 0x0AF0
		x"00",x"00",x"00",x"00",x"C0",x"C0",x"FE",x"FE", -- 0x0AF8
		x"FF",x"FF",x"FF",x"FF",x"F3",x"E3",x"E3",x"E3", -- 0x0B00
		x"E3",x"E3",x"C0",x"80",x"80",x"80",x"FF",x"FF", -- 0x0B08
		x"FE",x"FE",x"FC",x"FC",x"FC",x"FC",x"F0",x"E0", -- 0x0B10
		x"E0",x"E0",x"00",x"00",x"00",x"00",x"FE",x"FE", -- 0x0B18
		x"00",x"38",x"3B",x"3B",x"3B",x"3B",x"03",x"00", -- 0x0B20
		x"00",x"3E",x"3E",x"3E",x"3E",x"00",x"00",x"00", -- 0x0B28
		x"00",x"1E",x"9E",x"9E",x"80",x"9E",x"9E",x"1E", -- 0x0B30
		x"00",x"1E",x"1E",x"1E",x"00",x"00",x"00",x"00", -- 0x0B38
		x"00",x"33",x"33",x"33",x"03",x"00",x"3F",x"3F", -- 0x0B40
		x"3F",x"00",x"00",x"0E",x"0E",x"0E",x"0E",x"00", -- 0x0B48
		x"00",x"9E",x"9E",x"9E",x"80",x"00",x"00",x"78", -- 0x0B50
		x"78",x"78",x"00",x"EE",x"EE",x"EE",x"E0",x"00", -- 0x0B58
		x"00",x"1E",x"1E",x"1E",x"00",x"1E",x"1E",x"1E", -- 0x0B60
		x"00",x"00",x"00",x"0F",x"0F",x"0F",x"00",x"00", -- 0x0B68
		x"00",x"70",x"70",x"70",x"76",x"76",x"76",x"76", -- 0x0B70
		x"06",x"00",x"1C",x"9C",x"9C",x"80",x"00",x"00", -- 0x0B78
		x"00",x"3C",x"3C",x"3C",x"00",x"03",x"04",x"06", -- 0x0B80
		x"07",x"03",x"00",x"00",x"3C",x"3C",x"00",x"00", -- 0x0B88
		x"00",x"0C",x"12",x"1A",x"1E",x"0C",x"80",x"80", -- 0x0B90
		x"80",x"18",x"24",x"34",x"3C",x"18",x"00",x"00", -- 0x0B98
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA8
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC8
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0BD0
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0BD8
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BE8
		x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0BF0
		x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE", -- 0x0BF8
		x"A0",x"41",x"08",x"A9",x"97",x"E0",x"50",x"A9", -- 0x0C00
		x"B1",x"D8",x"5C",x"66",x"3B",x"BA",x"95",x"96", -- 0x0C08
		x"A0",x"98",x"D4",x"C0",x"A0",x"C2",x"28",x"14", -- 0x0C10
		x"00",x"88",x"88",x"24",x"95",x"0A",x"00",x"D8", -- 0x0C18
		x"CD",x"CD",x"86",x"83",x"99",x"6C",x"03",x"06", -- 0x0C20
		x"08",x"30",x"C0",x"21",x"57",x"89",x"71",x"8C", -- 0x0C28
		x"88",x"C4",x"A4",x"52",x"BD",x"D6",x"68",x"6A", -- 0x0C30
		x"6D",x"D0",x"CB",x"B5",x"52",x"40",x"A6",x"A4", -- 0x0C38
		x"C9",x"FC",x"4C",x"01",x"84",x"04",x"06",x"0C", -- 0x0C40
		x"18",x"B1",x"C7",x"9F",x"3F",x"C3",x"20",x"98", -- 0x0C48
		x"A8",x"C4",x"84",x"BA",x"DD",x"D6",x"68",x"6E", -- 0x0C50
		x"DD",x"66",x"36",x"B2",x"9B",x"1A",x"99",x"0D", -- 0x0C58
		x"C0",x"60",x"B2",x"5D",x"A2",x"9F",x"E9",x"60", -- 0x0C60
		x"06",x"1D",x"1D",x"8B",x"4F",x"4E",x"7C",x"90", -- 0x0C68
		x"08",x"54",x"24",x"1A",x"AD",x"3A",x"78",x"A5", -- 0x0C70
		x"5B",x"2D",x"86",x"90",x"39",x"7C",x"78",x"FB", -- 0x0C78
		x"80",x"10",x"21",x"23",x"3F",x"73",x"F0",x"81", -- 0x0C80
		x"86",x"08",x"90",x"A0",x"A0",x"40",x"C1",x"87", -- 0x0C88
		x"71",x"E3",x"C3",x"87",x"03",x"07",x"4E",x"9C", -- 0x0C90
		x"1C",x"1D",x"38",x"30",x"30",x"61",x"C1",x"37", -- 0x0C98
		x"7C",x"C8",x"01",x"33",x"CE",x"31",x"9C",x"CF", -- 0x0CA0
		x"71",x"1E",x"07",x"00",x"C0",x"E3",x"FF",x"FF", -- 0x0CA8
		x"BE",x"9C",x"00",x"01",x"61",x"73",x"BE",x"CC", -- 0x0CB0
		x"E0",x"1C",x"CF",x"20",x"1B",x"86",x"E0",x"FF", -- 0x0CB8
		x"FE",x"FC",x"FE",x"FC",x"FC",x"FE",x"FF",x"FF", -- 0x0CC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F3",x"C1",x"E5", -- 0x0CC8
		x"68",x"74",x"64",x"7A",x"3D",x"96",x"88",x"CE", -- 0x0CD0
		x"8D",x"C6",x"D6",x"E2",x"E3",x"73",x"19",x"35", -- 0x0CD8
		x"17",x"8B",x"CB",x"CA",x"C5",x"65",x"A4",x"D2", -- 0x0CE0
		x"12",x"09",x"09",x"89",x"E4",x"24",x"14",x"0A", -- 0x0CE8
		x"38",x"BC",x"54",x"52",x"50",x"A1",x"A1",x"52", -- 0x0CF0
		x"51",x"51",x"29",x"14",x"94",x"94",x"8A",x"4A", -- 0x0CF8
		x"82",x"82",x"C1",x"41",x"62",x"22",x"32",x"91", -- 0x0D00
		x"99",x"48",x"6C",x"04",x"06",x"82",x"43",x"61", -- 0x0D08
		x"04",x"05",x"0B",x"1A",x"32",x"34",x"18",x"08", -- 0x0D10
		x"09",x"89",x"8C",x"C4",x"45",x"43",x"22",x"22", -- 0x0D18
		x"71",x"38",x"18",x"0D",x"07",x"46",x"E0",x"F1", -- 0x0D20
		x"40",x"B3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D28
		x"E9",x"F2",x"CD",x"03",x"03",x"01",x"01",x"03", -- 0x0D30
		x"02",x"0A",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D38
		x"BE",x"BF",x"FE",x"ED",x"DF",x"FF",x"7F",x"FF", -- 0x0D40
		x"FF",x"EF",x"B7",x"FF",x"FF",x"FF",x"FF",x"DE", -- 0x0D48
		x"F7",x"FB",x"FB",x"8F",x"AF",x"79",x"3C",x"B6", -- 0x0D50
		x"C4",x"DF",x"F7",x"FF",x"FF",x"F5",x"21",x"33", -- 0x0D58
		x"54",x"4C",x"AA",x"A5",x"D3",x"CA",x"65",x"65", -- 0x0D60
		x"3C",x"1E",x"9E",x"49",x"4C",x"4C",x"22",x"21", -- 0x0D68
		x"3B",x"79",x"7C",x"72",x"32",x"99",x"4D",x"28", -- 0x0D70
		x"AC",x"A6",x"57",x"49",x"B6",x"B3",x"59",x"59", -- 0x0D78
		x"98",x"F6",x"DB",x"B7",x"41",x"31",x"0F",x"9B", -- 0x0D80
		x"F1",x"1C",x"CF",x"F8",x"61",x"06",x"8C",x"F8", -- 0x0D88
		x"48",x"A4",x"A4",x"A8",x"74",x"72",x"BA",x"D9", -- 0x0D90
		x"CC",x"27",x"D7",x"8B",x"C9",x"F4",x"7A",x"3A", -- 0x0D98
		x"07",x"00",x"C3",x"FF",x"4C",x"04",x"C0",x"E7", -- 0x0DA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DA8
		x"0E",x"E3",x"F0",x"30",x"1C",x"0F",x"C1",x"B8", -- 0x0DB0
		x"CE",x"E3",x"F1",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB8
		x"FF",x"7B",x"EF",x"FE",x"FF",x"FF",x"BF",x"FF", -- 0x0DC0
		x"FE",x"FE",x"7C",x"FC",x"FC",x"F8",x"F9",x"FC", -- 0x0DC8
		x"6F",x"FF",x"FC",x"EC",x"C8",x"8C",x"9E",x"5E", -- 0x0DD0
		x"4F",x"E7",x"F3",x"51",x"6D",x"24",x"16",x"93", -- 0x0DD8
		x"FE",x"F9",x"F0",x"F0",x"E0",x"F0",x"FD",x"E2", -- 0x0DE0
		x"F2",x"F9",x"D8",x"EC",x"E6",x"F1",x"D0",x"EC", -- 0x0DE8
		x"3F",x"07",x"81",x"C0",x"F0",x"7C",x"0E",x"E5", -- 0x0DF0
		x"73",x"3F",x"87",x"E1",x"30",x"0C",x"C7",x"70", -- 0x0DF8
		x"E6",x"F3",x"B8",x"E6",x"FB",x"FF",x"FF",x"FF", -- 0x0E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E08
		x"38",x"0F",x"85",x"E0",x"F8",x"FE",x"FF",x"FF", -- 0x0E10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E18
		x"FF",x"FF",x"FB",x"FF",x"FF",x"BD",x"FF",x"FF", -- 0x0E20
		x"FF",x"FF",x"FB",x"FF",x"BF",x"FF",x"FF",x"F7", -- 0x0E28
		x"FF",x"EF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF", -- 0x0E30
		x"FF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E38
		x"DF",x"FE",x"FF",x"FD",x"EF",x"FF",x"FF",x"FF", -- 0x0E40
		x"FF",x"FF",x"F7",x"BF",x"FB",x"FF",x"FF",x"FF", -- 0x0E48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E58
		x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"0E", -- 0x0E60
		x"2C",x"5C",x"4E",x"0F",x"87",x"C7",x"FF",x"FF", -- 0x0E68
		x"FF",x"7F",x"3F",x"03",x"4B",x"17",x"93",x"03", -- 0x0E70
		x"63",x"33",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E78
		x"FF",x"E7",x"E3",x"E0",x"F4",x"F1",x"F9",x"E0", -- 0x0E80
		x"C6",x"C3",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E88
		x"FF",x"FF",x"FF",x"3F",x"BF",x"79",x"38",x"38", -- 0x0E90
		x"1D",x"1C",x"FE",x"F8",x"F1",x"F0",x"F9",x"FF", -- 0x0E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EA0
		x"FF",x"7F",x"7F",x"AB",x"14",x"57",x"E8",x"1A", -- 0x0EA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EB0
		x"FF",x"FF",x"FF",x"7F",x"9F",x"66",x"C9",x"92", -- 0x0EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF", -- 0x0EC0
		x"0D",x"82",x"7A",x"AA",x"94",x"57",x"68",x"9A", -- 0x0EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0ED0
		x"FF",x"5F",x"94",x"69",x"BA",x"66",x"C9",x"92", -- 0x0ED8
		x"FF",x"FF",x"FF",x"FF",x"59",x"66",x"93",x"49", -- 0x0EE0
		x"AA",x"55",x"E6",x"4A",x"AD",x"B6",x"58",x"65", -- 0x0EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"17",x"18", -- 0x0EF0
		x"A4",x"4A",x"60",x"B7",x"45",x"9A",x"EC",x"69", -- 0x0EF8
		x"FF",x"57",x"B2",x"AE",x"D9",x"D7",x"7B",x"4B", -- 0x0F00
		x"FA",x"6F",x"FC",x"35",x"57",x"AA",x"6B",x"9A", -- 0x0F08
		x"FF",x"FF",x"FF",x"9D",x"67",x"DA",x"7F",x"64", -- 0x0F10
		x"DA",x"77",x"AA",x"D7",x"5A",x"AD",x"57",x"EC", -- 0x0F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"BB", -- 0x0F28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EA",x"D5",x"AA", -- 0x0F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F70
		x"FF",x"FD",x"F9",x"4A",x"F5",x"65",x"9A",x"AB", -- 0x0F78
		x"AF",x"9F",x"4F",x"7F",x"DF",x"7F",x"EF",x"5F", -- 0x0F80
		x"AF",x"7F",x"5F",x"AF",x"6F",x"9F",x"DF",x"6F", -- 0x0F88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"9E",x"43",x"49", -- 0x0FA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"59", -- 0x0FB8
		x"BF",x"7F",x"FF",x"4F",x"AD",x"B6",x"58",x"65", -- 0x0FC0
		x"95",x"6A",x"2D",x"96",x"59",x"66",x"93",x"49", -- 0x0FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"6B", -- 0x0FD0
		x"97",x"A9",x"2E",x"D5",x"29",x"EA",x"16",x"59", -- 0x0FD8
		x"5F",x"9F",x"7F",x"5F",x"9F",x"27",x"6F",x"97", -- 0x0FE0
		x"67",x"59",x"B6",x"AD",x"4A",x"E6",x"55",x"AA", -- 0x0FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF0
		x"FF",x"FF",x"DF",x"77",x"BF",x"66",x"5A",x"A5", -- 0x0FF8
		x"7F",x"3F",x"1F",x"0F",x"83",x"C1",x"C1",x"63", -- 0x1000
		x"6F",x"27",x"F7",x"B5",x"99",x"99",x"48",x"A5", -- 0x1008
		x"FF",x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x1010
		x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1018
		x"35",x"13",x"1D",x"09",x"0D",x"1D",x"3F",x"39", -- 0x1020
		x"7B",x"B3",x"A3",x"C3",x"C1",x"E1",x"E3",x"F7", -- 0x1028
		x"FF",x"7F",x"7F",x"BF",x"AF",x"8F",x"CF",x"CF", -- 0x1030
		x"87",x"87",x"CF",x"DF",x"DB",x"D3",x"C1",x"E1", -- 0x1038
		x"B1",x"75",x"B4",x"90",x"D9",x"9A",x"9C",x"C8", -- 0x1040
		x"68",x"58",x"6C",x"6C",x"6D",x"34",x"36",x"32", -- 0x1048
		x"EF",x"EF",x"EF",x"EF",x"E9",x"F1",x"71",x"33", -- 0x1050
		x"37",x"37",x"35",x"F8",x"F8",x"79",x"3B",x"3B", -- 0x1058
		x"FF",x"5F",x"8F",x"8F",x"CF",x"D7",x"E3",x"73", -- 0x1060
		x"77",x"35",x"39",x"39",x"1B",x"1C",x"0C",x"84", -- 0x1068
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"FF", -- 0x1070
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x1078
		x"86",x"C7",x"C7",x"C3",x"C3",x"E3",x"EF",x"61", -- 0x1080
		x"71",x"71",x"73",x"34",x"38",x"3B",x"1B",x"18", -- 0x1088
		x"3F",x"1F",x"7F",x"AF",x"AF",x"87",x"C7",x"C7", -- 0x1090
		x"9F",x"BF",x"D7",x"C3",x"A3",x"83",x"87",x"87", -- 0x1098
		x"65",x"2D",x"1D",x"16",x"0E",x"0A",x"1D",x"B6", -- 0x10A0
		x"D2",x"C3",x"C1",x"C1",x"E3",x"E3",x"66",x"2C", -- 0x10A8
		x"C3",x"E3",x"EF",x"DF",x"47",x"43",x"C3",x"C3", -- 0x10B0
		x"E7",x"2F",x"2F",x"6B",x"61",x"71",x"99",x"9B", -- 0x10B8
		x"90",x"98",x"8C",x"CC",x"55",x"2E",x"32",x"17", -- 0x10C0
		x"99",x"CB",x"DC",x"6C",x"26",x"23",x"15",x"17", -- 0x10C8
		x"6D",x"3E",x"77",x"B7",x"9F",x"1B",x"3B",x"7B", -- 0x10D0
		x"6C",x"9F",x"A7",x"63",x"A1",x"11",x"91",x"D8", -- 0x10D8
		x"BC",x"BE",x"51",x"21",x"30",x"78",x"78",x"7C", -- 0x10E0
		x"BD",x"DE",x"D6",x"E3",x"E1",x"E1",x"F0",x"F9", -- 0x10E8
		x"E0",x"60",x"78",x"3D",x"FD",x"9D",x"7E",x"CF", -- 0x10F0
		x"FF",x"EB",x"FF",x"79",x"6D",x"87",x"C7",x"E3", -- 0x10F8
		x"38",x"19",x"1E",x"1C",x"8E",x"CF",x"C7",x"E3", -- 0x1100
		x"61",x"71",x"38",x"18",x"18",x"58",x"CC",x"8C", -- 0x1108
		x"E1",x"70",x"30",x"18",x"18",x"38",x"F8",x"D8", -- 0x1110
		x"0C",x"8C",x"8C",x"84",x"44",x"5C",x"7C",x"7E", -- 0x1118
		x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1120
		x"FC",x"F8",x"E0",x"C0",x"E1",x"F3",x"E7",x"EF", -- 0x1128
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1130
		x"1F",x"0F",x"07",x"03",x"F3",x"F1",x"F8",x"FC", -- 0x1138
		x"F3",x"E3",x"E1",x"71",x"31",x"39",x"98",x"9C", -- 0x1140
		x"48",x"03",x"7F",x"FF",x"FF",x"FF",x"F9",x"F8", -- 0x1148
		x"FF",x"FF",x"DF",x"CF",x"C3",x"C1",x"C1",x"00", -- 0x1150
		x"E0",x"F0",x"F0",x"FC",x"FC",x"FE",x"9F",x"CF", -- 0x1158
		x"E0",x"67",x"9F",x"3F",x"FF",x"FF",x"FE",x"F8", -- 0x1160
		x"FC",x"F9",x"F7",x"EF",x"DF",x"BF",x"7F",x"7F", -- 0x1168
		x"07",x"C1",x"F1",x"F8",x"FC",x"FC",x"0E",x"07", -- 0x1170
		x"E3",x"F1",x"F9",x"FC",x"EC",x"E2",x"F0",x"F0", -- 0x1178
		x"FF",x"3F",x"9C",x"99",x"C3",x"C7",x"E7",x"CF", -- 0x1180
		x"9F",x"38",x"60",x"68",x"DB",x"B7",x"6F",x"6F", -- 0x1188
		x"F0",x"C0",x"00",x"78",x"FE",x"FF",x"FF",x"8F", -- 0x1190
		x"07",x"03",x"31",x"FC",x"FC",x"FE",x"FF",x"CF", -- 0x1198
		x"1E",x"6C",x"D9",x"B7",x"2F",x"5F",x"DF",x"FE", -- 0x11A0
		x"BD",x"37",x"6F",x"EF",x"DF",x"B3",x"61",x"40", -- 0x11A8
		x"01",x"F8",x"FE",x"FA",x"C0",x"98",x"7C",x"FF", -- 0x11B0
		x"FF",x"E3",x"00",x"00",x"80",x"98",x"3E",x"7F", -- 0x11B8
		x"20",x"20",x"71",x"79",x"73",x"37",x"17",x"07", -- 0x11C0
		x"05",x"0F",x"0B",x"03",x"01",x"80",x"80",x"8C", -- 0x11C8
		x"FF",x"F8",x"F8",x"FC",x"CE",x"C6",x"16",x"0C", -- 0x11D0
		x"81",x"C7",x"CF",x"9F",x"BF",x"3F",x"7F",x"7F", -- 0x11D8
		x"8E",x"0F",x"06",x"02",x"10",x"39",x"39",x"3A", -- 0x11E0
		x"38",x"38",x"30",x"00",x"0C",x"10",x"30",x"01", -- 0x11E8
		x"7C",x"70",x"EC",x"DC",x"D8",x"93",x"07",x"07", -- 0x11F0
		x"06",x"CC",x"CE",x"5B",x"11",x"20",x"2E",x"8D", -- 0x11F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"FC",x"F8", -- 0x1200
		x"F0",x"F9",x"FC",x"DC",x"8A",x"04",x"14",x"88", -- 0x1208
		x"F1",x"E1",x"C2",x"8D",x"C2",x"C8",x"30",x"A0", -- 0x1210
		x"48",x"58",x"0C",x"06",x"02",x"45",x"23",x"13", -- 0x1218
		x"81",x"03",x"07",x"0F",x"03",x"01",x"00",x"00", -- 0x1220
		x"00",x"18",x"0C",x"66",x"62",x"60",x"E0",x"20", -- 0x1228
		x"93",x"CD",x"DB",x"B7",x"AF",x"62",x"C1",x"8B", -- 0x1230
		x"1B",x"0B",x"07",x"17",x"1F",x"0E",x"0E",x"0C", -- 0x1238
		x"00",x"08",x"00",x"00",x"11",x"10",x"00",x"00", -- 0x1240
		x"00",x"00",x"01",x"00",x"00",x"10",x"00",x"00", -- 0x1248
		x"0D",x"09",x"1B",x"93",x"B7",x"67",x"67",x"4F", -- 0x1250
		x"0F",x"9F",x"1F",x"0F",x"06",x"00",x"00",x"00", -- 0x1258
		x"00",x"30",x"00",x"00",x"70",x"D0",x"30",x"21", -- 0x1260
		x"A0",x"A2",x"43",x"43",x"27",x"21",x"30",x"10", -- 0x1268
		x"80",x"40",x"70",x"39",x"19",x"01",x"00",x"00", -- 0x1270
		x"C0",x"30",x"86",x"E6",x"E0",x"C0",x"0C",x"18", -- 0x1278
		x"66",x"60",x"20",x"18",x"0C",x"06",x"02",x"00", -- 0x1280
		x"60",x"70",x"70",x"70",x"70",x"30",x"09",x"61", -- 0x1288
		x"05",x"1B",x"02",x"21",x"25",x"1D",x"28",x"48", -- 0x1290
		x"00",x"60",x"90",x"91",x"63",x"C3",x"23",x"21", -- 0x1298
		x"70",x"30",x"00",x"24",x"08",x"01",x"80",x"C0", -- 0x12A0
		x"80",x"80",x"00",x"48",x"01",x"44",x"E2",x"E4", -- 0x12A8
		x"00",x"06",x"0F",x"4F",x"9F",x"1F",x"06",x"00", -- 0x12B0
		x"1E",x"9E",x"CA",x"80",x"86",x"02",x"40",x"08", -- 0x12B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12D0
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12D8
		x"FF",x"FF",x"EF",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x12E0
		x"FF",x"BF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF", -- 0x12E8
		x"F9",x"F4",x"FA",x"F9",x"FC",x"FE",x"CF",x"C6", -- 0x12F0
		x"C0",x"A4",x"08",x"C0",x"E0",x"F0",x"F0",x"30", -- 0x12F8
		x"FF",x"FE",x"FE",x"FE",x"FE",x"FC",x"FF",x"FF", -- 0x1300
		x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FE", -- 0x1308
		x"10",x"00",x"00",x"00",x"00",x"80",x"03",x"C3", -- 0x1310
		x"C7",x"07",x"01",x"00",x"00",x"07",x"07",x"07", -- 0x1318
		x"FC",x"FF",x"FF",x"FD",x"F8",x"F8",x"F8",x"F8", -- 0x1320
		x"F8",x"FC",x"F4",x"F0",x"F0",x"F8",x"E4",x"E0", -- 0x1328
		x"00",x"00",x"80",x"80",x"90",x"18",x"00",x"00", -- 0x1330
		x"00",x"01",x"70",x"00",x"00",x"40",x"20",x"00", -- 0x1338
		x"F0",x"F0",x"F8",x"E8",x"C0",x"E0",x"F0",x"F8", -- 0x1340
		x"F8",x"F8",x"F4",x"C0",x"C0",x"E0",x"C8",x"C6", -- 0x1348
		x"04",x"04",x"4C",x"6C",x"28",x"18",x"D8",x"D8", -- 0x1350
		x"D8",x"D8",x"D8",x"2C",x"2C",x"6C",x"76",x"06", -- 0x1358
		x"E0",x"F0",x"F8",x"DC",x"C0",x"F0",x"F8",x"F8", -- 0x1360
		x"F8",x"C0",x"E0",x"E4",x"EC",x"E0",x"FC",x"EC", -- 0x1368
		x"36",x"34",x"00",x"20",x"30",x"71",x"01",x"03", -- 0x1370
		x"33",x"63",x"81",x"20",x"80",x"E0",x"80",x"30", -- 0x1378
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1380
		x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1388
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1390
		x"FF",x"7F",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1398
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF", -- 0x13A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13F8
		x"B6",x"76",x"F5",x"E4",x"EC",x"6C",x"CA",x"EB", -- 0x1400
		x"F9",x"98",x"98",x"D8",x"F6",x"B7",x"37",x"F7", -- 0x1408
		x"F8",x"F8",x"F8",x"FE",x"7F",x"33",x"31",x"31", -- 0x1410
		x"F1",x"FD",x"FF",x"EF",x"E7",x"E3",x"E1",x"E1", -- 0x1418
		x"F0",x"F9",x"FD",x"CD",x"C7",x"83",x"83",x"01", -- 0x1420
		x"01",x"0D",x"0D",x"0D",x"09",x"9F",x"F7",x"FD", -- 0x1428
		x"F8",x"CF",x"C7",x"C3",x"C3",x"C7",x"B7",x"BF", -- 0x1430
		x"DF",x"DF",x"8F",x"8F",x"9F",x"7F",x"7F",x"FF", -- 0x1438
		x"A5",x"48",x"99",x"9B",x"B7",x"FF",x"23",x"63", -- 0x1440
		x"63",x"C7",x"C7",x"A7",x"7F",x"FF",x"FF",x"FF", -- 0x1448
		x"FF",x"FF",x"FF",x"FF",x"FB",x"FF",x"FF",x"FF", -- 0x1450
		x"FF",x"FF",x"FF",x"EF",x"F7",x"FF",x"FF",x"FF", -- 0x1458
		x"0D",x"0F",x"99",x"98",x"38",x"FA",x"F7",x"E1", -- 0x1460
		x"EB",x"DF",x"DF",x"8E",x"1C",x"9D",x"98",x"BC", -- 0x1468
		x"66",x"C5",x"C5",x"C5",x"84",x"8C",x"BC",x"3C", -- 0x1470
		x"38",x"18",x"18",x"D8",x"FA",x"F3",x"F7",x"E7", -- 0x1478
		x"F8",x"FF",x"FF",x"FF",x"FF",x"FE",x"FD",x"DD", -- 0x1480
		x"DF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF", -- 0x1488
		x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1490
		x"FF",x"DE",x"9C",x"98",x"3A",x"7B",x"F7",x"F7", -- 0x1498
		x"F8",x"30",x"65",x"6F",x"67",x"C6",x"C6",x"8C", -- 0x14A0
		x"0C",x"18",x"1A",x"33",x"27",x"47",x"86",x"8C", -- 0x14A8
		x"EF",x"CF",x"87",x"0C",x"19",x"3B",x"23",x"6F", -- 0x14B0
		x"4F",x"5E",x"9C",x"BC",x"3C",x"78",x"62",x"E6", -- 0x14B8
		x"1B",x"39",x"31",x"71",x"E5",x"EF",x"CF",x"CE", -- 0x14C0
		x"8E",x"06",x"8C",x"8A",x"DA",x"F4",x"74",x"6C", -- 0x14C8
		x"CC",x"9C",x"98",x"18",x"19",x"39",x"71",x"F1", -- 0x14D0
		x"71",x"61",x"67",x"77",x"F7",x"F3",x"E3",x"6F", -- 0x14D8
		x"1B",x"79",x"79",x"FB",x"F3",x"F3",x"F1",x"F1", -- 0x14E0
		x"E1",x"E3",x"E3",x"C3",x"C7",x"C7",x"CF",x"BE", -- 0x14E8
		x"E7",x"D7",x"DB",x"DF",x"DF",x"CF",x"87",x"87", -- 0x14F0
		x"C7",x"D7",x"BF",x"9F",x"9F",x"1F",x"1F",x"BF", -- 0x14F8
		x"BD",x"7D",x"FC",x"F9",x"F9",x"F9",x"F3",x"F3", -- 0x1500
		x"F3",x"EF",x"CF",x"CF",x"8F",x"BF",x"3F",x"3F", -- 0x1508
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1510
		x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1518
		x"01",x"11",x"10",x"18",x"08",x"38",x"38",x"38", -- 0x1520
		x"38",x"38",x"30",x"00",x"06",x"1E",x"0F",x"0E", -- 0x1528
		x"CE",x"CF",x"07",x"47",x"C7",x"C3",x"81",x"61", -- 0x1530
		x"74",x"27",x"13",x"18",x"1C",x"0C",x"00",x"01", -- 0x1538
		x"8C",x"88",x"C0",x"C1",x"C3",x"C3",x"C3",x"81", -- 0x1540
		x"01",x"10",x"30",x"70",x"78",x"70",x"20",x"26", -- 0x1548
		x"00",x"01",x"01",x"B3",x"9F",x"CF",x"E7",x"F1", -- 0x1550
		x"EC",x"D6",x"07",x"0F",x"1E",x"0F",x"03",x"03", -- 0x1558
		x"0C",x"09",x"83",x"C7",x"E3",x"60",x"30",x"8C", -- 0x1560
		x"C6",x"C3",x"41",x"A0",x"B0",x"98",x"4C",x"20", -- 0x1568
		x"07",x"26",x"98",x"E2",x"FE",x"FF",x"3D",x"03", -- 0x1570
		x"0F",x"0C",x"9B",x"C1",x"78",x"00",x"08",x"01", -- 0x1578
		x"60",x"60",x"34",x"1B",x"0C",x"0F",x"03",x"80", -- 0x1580
		x"C0",x"E0",x"C0",x"C1",x"99",x"1C",x"3F",x"3F", -- 0x1588
		x"CF",x"1F",x"3E",x"FC",x"FC",x"31",x"83",x"F7", -- 0x1590
		x"6F",x"1F",x"7F",x"FF",x"FF",x"78",x"00",x"F0", -- 0x1598
		x"BF",x"9F",x"83",x"C0",x"60",x"70",x"39",x"1E", -- 0x15A0
		x"07",x"01",x"00",x"80",x"03",x"9F",x"07",x"00", -- 0x15A8
		x"F0",x"F0",x"E2",x"6C",x"1C",x"F8",x"F0",x"E2", -- 0x15B0
		x"0E",x"FE",x"1C",x"7C",x"F8",x"F1",x"C1",x"33", -- 0x15B8
		x"31",x"03",x"00",x"00",x"01",x"07",x"03",x"48", -- 0x15C0
		x"DC",x"98",x"B9",x"B1",x"71",x"61",x"83",x"C3", -- 0x15C8
		x"8F",x"1F",x"3E",x"FC",x"FC",x"F0",x"F0",x"E0", -- 0x15D0
		x"00",x"C1",x"C1",x"C3",x"C7",x"EF",x"CF",x"9F", -- 0x15D8
		x"E0",x"E0",x"F1",x"F9",x"FC",x"FF",x"FF",x"FF", -- 0x15E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E8
		x"1C",x"78",x"F1",x"E3",x"03",x"E7",x"EF",x"FF", -- 0x15F0
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"FF",x"FF", -- 0x15F8
		x"E4",x"80",x"49",x"09",x"80",x"00",x"80",x"C0", -- 0x1600
		x"C9",x"C9",x"C8",x"C8",x"84",x"02",x"21",x"70", -- 0x1608
		x"8E",x"02",x"81",x"87",x"80",x"80",x"08",x"1E", -- 0x1610
		x"1E",x"1E",x"1E",x"1C",x"00",x"03",x"87",x"84", -- 0x1618
		x"61",x"09",x"31",x"70",x"70",x"70",x"78",x"60", -- 0x1620
		x"00",x"02",x"06",x"0C",x"19",x"21",x"60",x"66", -- 0x1628
		x"21",x"23",x"A3",x"A3",x"91",x"91",x"C0",x"40", -- 0x1630
		x"48",x"08",x"08",x"24",x"20",x"12",x"13",x"01", -- 0x1638
		x"F0",x"F0",x"E1",x"E7",x"C3",x"C3",x"E2",x"E0", -- 0x1640
		x"E1",x"F1",x"10",x"30",x"70",x"30",x"39",x"1B", -- 0x1648
		x"9C",x"8E",x"C0",x"C0",x"E3",x"A7",x"32",x"F0", -- 0x1650
		x"F0",x"B9",x"1F",x"3D",x"74",x"E4",x"C4",x"84", -- 0x1658
		x"13",x"12",x"10",x"08",x"00",x"06",x"00",x"10", -- 0x1660
		x"90",x"90",x"91",x"81",x"80",x"C8",x"C8",x"C4", -- 0x1668
		x"18",x"10",x"20",x"04",x"0F",x"1F",x"1F",x"0F", -- 0x1670
		x"0F",x"07",x"07",x"87",x"C3",x"43",x"01",x"01", -- 0x1678
		x"30",x"F0",x"72",x"7B",x"67",x"04",x"08",x"01", -- 0x1680
		x"01",x"03",x"0F",x"0F",x"0F",x"87",x"83",x"C1", -- 0x1688
		x"10",x"11",x"11",x"10",x"18",x"88",x"88",x"1C", -- 0x1690
		x"0C",x"02",x"83",x"C7",x"C7",x"E3",x"F1",x"BC", -- 0x1698
		x"80",x"00",x"00",x"80",x"D8",x"FC",x"F8",x"F0", -- 0x16A0
		x"F8",x"FC",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16A8
		x"18",x"38",x"70",x"60",x"06",x"0C",x"18",x"08", -- 0x16B0
		x"04",x"00",x"80",x"C0",x"8C",x"D2",x"F1",x"F9", -- 0x16B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF", -- 0x16C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16D8
		x"C2",x"E4",x"FC",x"FC",x"E4",x"E0",x"C0",x"F8", -- 0x16E0
		x"F8",x"F8",x"F8",x"F8",x"F8",x"E0",x"C0",x"C4", -- 0x16E8
		x"C0",x"C0",x"00",x"00",x"E1",x"E0",x"00",x"00", -- 0x16F0
		x"03",x"71",x"01",x"00",x"18",x"00",x"34",x"06", -- 0x16F8
		x"FC",x"FC",x"FC",x"E4",x"C0",x"C0",x"E8",x"F8", -- 0x1700
		x"F8",x"F8",x"F8",x"F8",x"C0",x"C0",x"E0",x"E0", -- 0x1708
		x"06",x"06",x"6C",x"0C",x"0C",x"D8",x"D8",x"D8", -- 0x1710
		x"D8",x"D8",x"18",x"08",x"6C",x"6C",x"04",x"04", -- 0x1718
		x"F4",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC", -- 0x1720
		x"F8",x"F8",x"FA",x"FC",x"F9",x"FF",x"FF",x"FC", -- 0x1728
		x"01",x"21",x"41",x"01",x"11",x"31",x"01",x"00", -- 0x1730
		x"00",x"08",x"18",x"90",x"80",x"80",x"00",x"00", -- 0x1738
		x"FE",x"F9",x"F8",x"FC",x"FE",x"FF",x"FF",x"FF", -- 0x1740
		x"FF",x"FC",x"FC",x"FC",x"FF",x"FE",x"FE",x"FE", -- 0x1748
		x"27",x"C7",x"87",x"00",x"00",x"81",x"87",x"87", -- 0x1750
		x"03",x"03",x"01",x"C1",x"81",x"01",x"01",x"20", -- 0x1758
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1760
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1768
		x"30",x"F0",x"F0",x"E0",x"C0",x"88",x"D8",x"FC", -- 0x1770
		x"FC",x"FE",x"FC",x"FD",x"F9",x"FB",x"F7",x"FF", -- 0x1778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x1780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1788
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1790
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17C0
		x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17D8
		x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x17E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F0
		x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F8
		x"FF",x"FE",x"FF",x"F7",x"F7",x"FE",x"FF",x"FF", -- 0x1800
		x"FF",x"FF",x"FF",x"DF",x"FF",x"FF",x"FE",x"FF", -- 0x1808
		x"76",x"0A",x"21",x"89",x"4B",x"01",x"80",x"43", -- 0x1810
		x"A0",x"C0",x"41",x"9C",x"EC",x"A6",x"D6",x"F3", -- 0x1818
		x"42",x"C1",x"21",x"81",x"46",x"43",x"91",x"11", -- 0x1820
		x"00",x"44",x"80",x"E0",x"D4",x"F5",x"BA",x"FF", -- 0x1828
		x"7E",x"0A",x"29",x"09",x"CB",x"01",x"C0",x"03", -- 0x1830
		x"21",x"01",x"40",x"1C",x"0A",x"45",x"D6",x"F3", -- 0x1838
		x"42",x"51",x"39",x"8D",x"42",x"D4",x"FA",x"DB", -- 0x1840
		x"E0",x"E0",x"C0",x"E8",x"F0",x"F8",x"B2",x"FE", -- 0x1848
		x"7E",x"0A",x"09",x"89",x"8B",x"01",x"80",x"13", -- 0x1850
		x"01",x"01",x"01",x"3F",x"25",x"20",x"20",x"F5", -- 0x1858
		x"68",x"40",x"00",x"00",x"81",x"80",x"81",x"01", -- 0x1860
		x"00",x"A1",x"D0",x"E0",x"EC",x"FA",x"FF",x"FE", -- 0x1868
		x"7E",x"08",x"09",x"08",x"8A",x"01",x"80",x"62", -- 0x1870
		x"20",x"01",x"41",x"5D",x"40",x"E0",x"D0",x"FD", -- 0x1878
		x"42",x"61",x"21",x"89",x"44",x"C1",x"90",x"EC", -- 0x1880
		x"F9",x"FE",x"BD",x"FF",x"FF",x"FF",x"F6",x"FF", -- 0x1888
		x"7E",x"0A",x"09",x"09",x"8B",x"01",x"80",x"83", -- 0x1890
		x"20",x"C5",x"2B",x"9F",x"FD",x"FF",x"EF",x"FF", -- 0x1898
		x"42",x"C1",x"21",x"83",x"47",x"47",x"93",x"05", -- 0x18A0
		x"83",x"47",x"0F",x"8F",x"0D",x"5F",x"3F",x"FF", -- 0x18A8
		x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD", -- 0x18B0
		x"FF",x"BF",x"FF",x"FF",x"EF",x"FB",x"FB",x"DF", -- 0x18B8
		x"82",x"24",x"46",x"A8",x"9C",x"50",x"40",x"24", -- 0x18C0
		x"B0",x"80",x"08",x"80",x"0A",x"07",x"37",x"BF", -- 0x18C8
		x"02",x"41",x"00",x"20",x"A0",x"01",x"50",x"2C", -- 0x18D0
		x"21",x"97",x"2F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x18D8
		x"42",x"C1",x"21",x"81",x"44",x"43",x"91",x"11", -- 0x18E0
		x"F0",x"54",x"00",x"98",x"08",x"50",x"0C",x"A0", -- 0x18E8
		x"7E",x"0B",x"09",x"01",x"0B",x"03",x"87",x"13", -- 0x18F0
		x"03",x"07",x"0D",x"7F",x"3F",x"3F",x"7B",x"FF", -- 0x18F8
		x"42",x"C1",x"21",x"81",x"44",x"42",x"91",x"10", -- 0x1900
		x"F2",x"5F",x"0F",x"8D",x"0F",x"5F",x"3F",x"FF", -- 0x1908
		x"7E",x"0B",x"09",x"09",x"8B",x"03",x"97",x"7D", -- 0x1910
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x1918
		x"42",x"C1",x"21",x"81",x"56",x"43",x"90",x"10", -- 0x1920
		x"3B",x"FF",x"BF",x"FF",x"FF",x"FF",x"EF",x"FF", -- 0x1928
		x"7E",x"0B",x"09",x"09",x"8B",x"03",x"97",x"BF", -- 0x1930
		x"FF",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1938
		x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1940
		x"DF",x"FF",x"FF",x"FF",x"FE",x"FD",x"FE",x"FE", -- 0x1948
		x"FA",x"E8",x"C4",x"E4",x"92",x"E0",x"C9",x"B4", -- 0x1950
		x"E2",x"95",x"46",x"8A",x"42",x"07",x"6B",x"4D", -- 0x1958
		x"FF",x"FF",x"FF",x"FD",x"F0",x"F8",x"E0",x"C4", -- 0x1960
		x"B0",x"80",x"0C",x"80",x"0D",x"23",x"34",x"93", -- 0x1968
		x"FE",x"FD",x"E8",x"B0",x"20",x"01",x"50",x"2C", -- 0x1970
		x"22",x"91",x"19",x"91",x"40",x"B1",x"49",x"33", -- 0x1978
		x"FF",x"FE",x"F8",x"FC",x"F4",x"F8",x"E0",x"EC", -- 0x1980
		x"F0",x"E4",x"D4",x"C8",x"8C",x"C3",x"54",x"F3", -- 0x1988
		x"02",x"01",x"40",x"40",x"A0",x"21",x"50",x"2C", -- 0x1990
		x"3A",x"91",x"19",x"91",x"40",x"31",x"49",x"33", -- 0x1998
		x"FF",x"DF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x19A0
		x"FD",x"FA",x"FC",x"FC",x"B8",x"B3",x"34",x"93", -- 0x19A8
		x"FD",x"FB",x"F2",x"D0",x"A0",x"81",x"50",x"8C", -- 0x19B0
		x"3A",x"91",x"19",x"91",x"40",x"31",x"49",x"33", -- 0x19B8
		x"FF",x"FF",x"BF",x"FF",x"FF",x"FB",x"FF",x"FF", -- 0x19C0
		x"FF",x"FE",x"FF",x"FC",x"FD",x"E3",x"34",x"90", -- 0x19C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF", -- 0x19D0
		x"FA",x"B1",x"45",x"A9",x"C2",x"87",x"6B",x"4D", -- 0x19D8
		x"2F",x"9F",x"07",x"8B",x"01",x"A1",x"04",x"04", -- 0x19E0
		x"D0",x"8C",x"0C",x"80",x"0D",x"22",x"35",x"90", -- 0x19E8
		x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x19F0
		x"FF",x"FF",x"F7",x"F7",x"7F",x"FF",x"FF",x"FF", -- 0x19F8
		x"7F",x"97",x"07",x"81",x"0C",x"A0",x"00",x"24", -- 0x1A00
		x"B0",x"84",x"08",x"80",x"0D",x"23",x"34",x"90", -- 0x1A08
		x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"7F",x"3F", -- 0x1A10
		x"19",x"90",x"54",x"A9",x"C2",x"87",x"6B",x"4D", -- 0x1A18
		x"A6",x"44",x"00",x"89",x"04",x"A0",x"00",x"24", -- 0x1A20
		x"B0",x"84",x"08",x"80",x"0D",x"23",x"34",x"90", -- 0x1A28
		x"FF",x"7F",x"7F",x"BF",x"BF",x"BF",x"77",x"33", -- 0x1A30
		x"23",x"93",x"57",x"23",x"81",x"81",x"69",x"4C", -- 0x1A38
		x"6F",x"9F",x"0F",x"8B",x"01",x"A1",x"00",x"05", -- 0x1A40
		x"D0",x"8C",x"0C",x"80",x"0D",x"22",x"34",x"90", -- 0x1A48
		x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"BF",x"7F", -- 0x1A50
		x"7F",x"FF",x"FF",x"EF",x"C3",x"87",x"6B",x"4D", -- 0x1A58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"B8", -- 0x1A60
		x"A0",x"80",x"08",x"84",x"01",x"2B",x"3C",x"90", -- 0x1A68
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F", -- 0x1A70
		x"7F",x"5F",x"17",x"03",x"C3",x"83",x"69",x"4C", -- 0x1A78
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F5", -- 0x1A80
		x"D0",x"54",x"00",x"90",x"08",x"50",x"0C",x"A0", -- 0x1A88
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"FF",x"67", -- 0x1A90
		x"00",x"00",x"00",x"26",x"05",x"20",x"20",x"C5", -- 0x1A98
		x"42",x"C1",x"21",x"81",x"44",x"40",x"90",x"14", -- 0x1AA0
		x"3D",x"FF",x"FE",x"FB",x"FF",x"FF",x"FF",x"FF", -- 0x1AA8
		x"7E",x"0A",x"81",x"09",x"8B",x"01",x"00",x"25", -- 0x1AB0
		x"00",x"80",x"41",x"97",x"FF",x"F7",x"FF",x"FF", -- 0x1AB8
		x"FE",x"FC",x"FE",x"FD",x"F8",x"FC",x"BE",x"FE", -- 0x1AC0
		x"FC",x"F8",x"FE",x"FC",x"FC",x"F8",x"FC",x"FE", -- 0x1AC8
		x"7E",x"0A",x"01",x"09",x"0B",x"01",x"00",x"13", -- 0x1AD0
		x"01",x"01",x"01",x"33",x"25",x"30",x"20",x"F5", -- 0x1AD8
		x"A4",x"40",x"06",x"89",x"0C",x"A0",x"00",x"44", -- 0x1AE0
		x"C0",x"80",x"08",x"81",x"00",x"22",x"35",x"90", -- 0x1AE8
		x"FF",x"7F",x"7F",x"7F",x"BF",x"3F",x"7F",x"3B", -- 0x1AF0
		x"7F",x"3F",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x1AF8
		x"BF",x"BB",x"FF",x"FA",x"DF",x"FF",x"FB",x"EF", -- 0x1B00
		x"EF",x"EF",x"FF",x"BF",x"BB",x"BB",x"FF",x"FF", -- 0x1B08
		x"7D",x"75",x"FF",x"DB",x"DB",x"7B",x"7F",x"DD", -- 0x1B10
		x"DD",x"7F",x"EF",x"EF",x"FF",x"FB",x"7B",x"7E", -- 0x1B18
		x"FF",x"FB",x"BB",x"FF",x"FF",x"FE",x"DC",x"DD", -- 0x1B20
		x"FD",x"FF",x"EF",x"ED",x"FF",x"FF",x"F7",x"FF", -- 0x1B28
		x"7F",x"FB",x"FB",x"DB",x"FF",x"FF",x"FF",x"DF", -- 0x1B30
		x"DF",x"F7",x"FF",x"FE",x"7E",x"7F",x"EF",x"EF", -- 0x1B38
		x"FF",x"FB",x"BB",x"FF",x"FF",x"FE",x"DC",x"DD", -- 0x1B40
		x"FD",x"FF",x"EF",x"ED",x"FF",x"FF",x"F7",x"FF", -- 0x1B48
		x"7C",x"FA",x"FB",x"DA",x"FF",x"FF",x"FF",x"DF", -- 0x1B50
		x"DF",x"F7",x"FF",x"FE",x"7E",x"7F",x"EF",x"EF", -- 0x1B58
		x"82",x"24",x"46",x"E8",x"BC",x"50",x"40",x"24", -- 0x1B60
		x"B0",x"8C",x"0C",x"80",x"0D",x"23",x"34",x"93", -- 0x1B68
		x"02",x"41",x"20",x"20",x"A0",x"21",x"50",x"2C", -- 0x1B70
		x"3A",x"91",x"19",x"91",x"40",x"B1",x"49",x"33", -- 0x1B78
		x"42",x"C1",x"21",x"81",x"46",x"43",x"91",x"11", -- 0x1B80
		x"F0",x"54",x"00",x"98",x"08",x"50",x"0C",x"A0", -- 0x1B88
		x"7E",x"0A",x"09",x"09",x"8B",x"01",x"80",x"13", -- 0x1B90
		x"01",x"01",x"01",x"3F",x"25",x"20",x"20",x"F5", -- 0x1B98
		x"A6",x"42",x"03",x"81",x"0C",x"A0",x"00",x"24", -- 0x1BA0
		x"B0",x"8C",x"0C",x"80",x"0D",x"23",x"34",x"90", -- 0x1BA8
		x"08",x"10",x"20",x"A4",x"A2",x"B0",x"5B",x"2E", -- 0x1BB0
		x"2A",x"99",x"55",x"A9",x"C2",x"87",x"6B",x"4D", -- 0x1BB8
		x"FF",x"FF",x"FF",x"FF",x"E7",x"E3",x"E0",x"F4", -- 0x1BC0
		x"F1",x"F9",x"E0",x"C6",x"C3",x"E7",x"FF",x"FF", -- 0x1BC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"BF", -- 0x1BD0
		x"7F",x"3F",x"3F",x"1F",x"1F",x"FF",x"FF",x"FF", -- 0x1BD8
		x"FF",x"FF",x"FF",x"FF",x"E7",x"E3",x"E0",x"F4", -- 0x1BE0
		x"F1",x"F9",x"E0",x"C6",x"C3",x"E7",x"FF",x"FF", -- 0x1BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"BF", -- 0x1BF0
		x"7F",x"3F",x"3F",x"1F",x"1F",x"FF",x"FF",x"FF", -- 0x1BF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"00", -- 0x1C08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"00",x"00", -- 0x1C18
		x"FF",x"FF",x"7B",x"42",x"FF",x"00",x"CF",x"FF", -- 0x1C20
		x"18",x"18",x"18",x"1C",x"1C",x"1C",x"1C",x"1C", -- 0x1C28
		x"FF",x"00",x"DF",x"13",x"FF",x"03",x"FC",x"FF", -- 0x1C30
		x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
		x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C", -- 0x1C40
		x"1C",x"FF",x"00",x"3E",x"41",x"00",x"00",x"00", -- 0x1C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
		x"07",x"FC",x"00",x"00",x"00",x"00",x"00",x"18", -- 0x1C58
		x"FF",x"FF",x"FF",x"00",x"00",x"2F",x"EF",x"FF", -- 0x1C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C68
		x"F2",x"E7",x"40",x"00",x"00",x"BE",x"BE",x"FF", -- 0x1C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C78
		x"FF",x"FE",x"8E",x"9C",x"9C",x"BF",x"5F",x"1F", -- 0x1C80
		x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C88
		x"2F",x"97",x"17",x"2F",x"FF",x"FF",x"FF",x"FF", -- 0x1C90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C98
		x"1F",x"07",x"FF",x"C3",x"7B",x"FB",x"7F",x"4F", -- 0x1CA0
		x"9F",x"BF",x"BF",x"BF",x"3E",x"3E",x"3E",x"29", -- 0x1CA8
		x"F8",x"FF",x"FF",x"FF",x"FF",x"BF",x"7F",x"FF", -- 0x1CB0
		x"FB",x"EF",x"1C",x"99",x"D3",x"42",x"06",x"C2", -- 0x1CB8
		x"2F",x"FF",x"02",x"2C",x"2F",x"20",x"3E",x"17", -- 0x1CC0
		x"09",x"84",x"C2",x"61",x"B0",x"B8",x"1C",x"4F", -- 0x1CC8
		x"D2",x"D2",x"92",x"52",x"D2",x"12",x"1B",x"09", -- 0x1CD0
		x"00",x"80",x"C0",x"60",x"30",x"00",x"00",x"00", -- 0x1CD8
		x"F9",x"00",x"00",x"00",x"FF",x"FF",x"02",x"7D", -- 0x1CE0
		x"7D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CE8
		x"FF",x"00",x"00",x"00",x"FF",x"F7",x"00",x"F7", -- 0x1CF0
		x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"41",x"01", -- 0x1D08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D18
		x"3F",x"E0",x"EC",x"CF",x"C9",x"CA",x"C8",x"C3", -- 0x1D20
		x"1E",x"60",x"80",x"40",x"20",x"00",x"00",x"00", -- 0x1D28
		x"FF",x"00",x"00",x"FF",x"FF",x"E0",x"1F",x"FF", -- 0x1D30
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
		x"00",x"00",x"00",x"00",x"20",x"C0",x"E0",x"3E", -- 0x1D40
		x"03",x"00",x"04",x"00",x"07",x"81",x"C0",x"E0", -- 0x1D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
		x"E0",x"3F",x"80",x"40",x"80",x"00",x"00",x"00", -- 0x1D58
		x"F8",x"38",x"38",x"00",x"00",x"00",x"EF",x"EF", -- 0x1D60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D68
		x"FF",x"81",x"81",x"81",x"00",x"00",x"BE",x"BE", -- 0x1D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D78
		x"A2",x"F2",x"E9",x"E0",x"C2",x"CF",x"FF",x"FF", -- 0x1D80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D88
		x"7F",x"FF",x"71",x"6B",x"E1",x"E8",x"FC",x"FA", -- 0x1D90
		x"F8",x"F0",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D98
		x"FD",x"F1",x"E3",x"E7",x"CF",x"CF",x"CC",x"C8", -- 0x1DA0
		x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7", -- 0x1DA8
		x"80",x"18",x"3F",x"13",x"03",x"F3",x"08",x"00", -- 0x1DB0
		x"10",x"1F",x"1F",x"0F",x"00",x"20",x"3E",x"37", -- 0x1DB8
		x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7", -- 0x1DC0
		x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C3",x"C3", -- 0x1DC8
		x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3B", -- 0x1DD0
		x"3B",x"39",x"29",x"2C",x"22",x"02",x"08",x"80", -- 0x1DD8
		x"E3",x"F1",x"F1",x"F8",x"F8",x"FC",x"FE",x"FF", -- 0x1DE0
		x"00",x"FF",x"7D",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE8
		x"C3",x"E0",x"F0",x"F8",x"FF",x"FF",x"FF",x"00", -- 0x1DF0
		x"7F",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"00",x"00", -- 0x1E08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"00",x"00", -- 0x1E18
		x"3F",x"DB",x"C0",x"C0",x"E7",x"F0",x"17",x"10", -- 0x1E20
		x"FF",x"10",x"33",x"E1",x"0E",x"1C",x"7C",x"74", -- 0x1E28
		x"FC",x"7F",x"1F",x"1B",x"63",x"00",x"68",x"04", -- 0x1E30
		x"F0",x"7F",x"FC",x"71",x"E3",x"43",x"42",x"02", -- 0x1E38
		x"75",x"75",x"75",x"75",x"71",x"3F",x"1E",x"86", -- 0x1E40
		x"C0",x"70",x"7C",x"0E",x"00",x"00",x"00",x"00", -- 0x1E48
		x"80",x"02",x"83",x"03",x"81",x"80",x"40",x"00", -- 0x1E50
		x"00",x"00",x"00",x"3F",x"2F",x"2F",x"2F",x"31", -- 0x1E58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"CF",x"DB", -- 0x1E60
		x"17",x"06",x"0C",x"10",x"00",x"00",x"00",x"00", -- 0x1E68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"DD",x"6B", -- 0x1E70
		x"08",x"04",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
		x"F7",x"27",x"0F",x"13",x"02",x"04",x"04",x"00", -- 0x1E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
		x"FF",x"FF",x"FF",x"BF",x"9F",x"3F",x"17",x"03", -- 0x1E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
		x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00", -- 0x1EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
		x"FF",x"FF",x"A7",x"07",x"0F",x"0E",x"05",x"0D", -- 0x1EB0
		x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
		x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00", -- 0x1EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
		x"FF",x"3F",x"EF",x"8F",x"1F",x"3F",x"2F",x"13", -- 0x1ED0
		x"3F",x"3F",x"0B",x"07",x"07",x"1F",x"0B",x"01", -- 0x1ED8
		x"FF",x"3F",x"6B",x"4F",x"02",x"00",x"01",x"00", -- 0x1EE0
		x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7", -- 0x1EF0
		x"EF",x"4F",x"1F",x"17",x"0F",x"0F",x"1B",x"11", -- 0x1EF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F00
		x"6F",x"37",x"0F",x"0D",x"18",x"01",x"21",x"00", -- 0x1F08
		x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"FF",x"FF", -- 0x1F10
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x1F18
		x"FF",x"7F",x"3F",x"63",x"47",x"0F",x"0D",x"01", -- 0x1F20
		x"07",x"0D",x"09",x"03",x"07",x"04",x"01",x"00", -- 0x1F28
		x"FF",x"FF",x"BD",x"3B",x"FF",x"FF",x"FF",x"FF", -- 0x1F30
		x"FF",x"FF",x"FF",x"FF",x"FB",x"FF",x"FF",x"7F", -- 0x1F38
		x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00", -- 0x1F40
		x"01",x"03",x"05",x"00",x"02",x"01",x"00",x"00", -- 0x1F48
		x"FF",x"7F",x"3F",x"9B",x"7F",x"FF",x"7F",x"FF", -- 0x1F50
		x"FF",x"FF",x"7F",x"7F",x"7B",x"BD",x"BF",x"FF", -- 0x1F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"DF", -- 0x1F60
		x"1B",x"0E",x"06",x"0C",x"08",x"00",x"00",x"00", -- 0x1F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F70
		x"FF",x"CF",x"CF",x"9F",x"1B",x"03",x"01",x"01", -- 0x1F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1FB8
		x"E0",x"00",x"00",x"00",x"80",x"40",x"00",x"BE", -- 0x1FC0
		x"BE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC8
		x"2D",x"21",x"3E",x"00",x"00",x"00",x"7B",x"FB", -- 0x1FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD8
		x"E3",x"D7",x"C2",x"D1",x"F9",x"F4",x"F0",x"E1", -- 0x1FE0
		x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE8
		x"FF",x"1F",x"3F",x"3F",x"7F",x"BF",x"3F",x"7F", -- 0x1FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x1FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
