-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_A2 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_A2 is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"DF",x"B7",x"AF",x"8E",x"88",x"56",x"8D",x"C6", -- 0x0000
		x"84",x"81",x"53",x"A2",x"91",x"C5",x"CE",x"DE", -- 0x0008
		x"B4",x"6E",x"35",x"8C",x"73",x"F6",x"7E",x"F7", -- 0x0010
		x"73",x"2E",x"0D",x"20",x"91",x"06",x"A9",x"CF", -- 0x0018
		x"AA",x"54",x"55",x"AA",x"AA",x"55",x"AD",x"EA", -- 0x0020
		x"74",x"9E",x"87",x"27",x"BB",x"11",x"85",x"5E", -- 0x0028
		x"B4",x"AE",x"4D",x"55",x"A3",x"AA",x"44",x"55", -- 0x0030
		x"9A",x"8A",x"25",x"55",x"66",x"AB",x"AB",x"D5", -- 0x0038
		x"EE",x"4F",x"9B",x"D5",x"B1",x"4A",x"02",x"8F", -- 0x0040
		x"EA",x"55",x"DD",x"3A",x"09",x"91",x"C2",x"6E", -- 0x0048
		x"74",x"6A",x"E9",x"F4",x"E3",x"68",x"34",x"95", -- 0x0050
		x"9A",x"CA",x"E5",x"75",x"4E",x"9D",x"3F",x"FF", -- 0x0058
		x"FF",x"DF",x"0D",x"54",x"89",x"60",x"7E",x"1F", -- 0x0060
		x"2A",x"84",x"43",x"A4",x"F3",x"ED",x"DE",x"E6", -- 0x0068
		x"5C",x"3E",x"ED",x"F5",x"A3",x"9A",x"54",x"F5", -- 0x0070
		x"7A",x"CA",x"E5",x"54",x"25",x"B9",x"D9",x"FD", -- 0x0078
		x"B3",x"46",x"05",x"10",x"D8",x"7D",x"67",x"2E", -- 0x0080
		x"84",x"C3",x"07",x"6F",x"4F",x"1E",x"1A",x"3B", -- 0x0088
		x"FF",x"FA",x"B5",x"74",x"93",x"A8",x"C4",x"D5", -- 0x0090
		x"FA",x"C2",x"A1",x"55",x"66",x"AB",x"AB",x"55", -- 0x0098
		x"36",x"7C",x"D5",x"EA",x"AA",x"7D",x"B9",x"7A", -- 0x00A0
		x"F4",x"AA",x"DB",x"73",x"4D",x"2C",x"1E",x"BF", -- 0x00A8
		x"B4",x"AA",x"45",x"55",x"A3",x"AA",x"44",x"55", -- 0x00B0
		x"9A",x"AA",x"25",x"55",x"62",x"AB",x"CB",x"55", -- 0x00B8
		x"CA",x"6C",x"75",x"3C",x"DE",x"3C",x"7C",x"DA", -- 0x00C0
		x"EC",x"B6",x"72",x"23",x"0D",x"1F",x"BC",x"EE", -- 0x00C8
		x"B4",x"AE",x"4D",x"54",x"83",x"88",x"44",x"55", -- 0x00D0
		x"9A",x"82",x"21",x"55",x"66",x"EB",x"A9",x"D5", -- 0x00D8
		x"EE",x"57",x"0F",x"0F",x"D4",x"AE",x"33",x"FF", -- 0x00E0
		x"4B",x"A6",x"F5",x"21",x"49",x"09",x"84",x"EE", -- 0x00E8
		x"F4",x"A8",x"C5",x"55",x"A3",x"EA",x"44",x"55", -- 0x00F0
		x"DA",x"8A",x"A5",x"55",x"22",x"8B",x"AB",x"D5", -- 0x00F8
		x"EF",x"47",x"17",x"57",x"FE",x"7C",x"3C",x"0A", -- 0x0100
		x"44",x"A6",x"72",x"73",x"5F",x"AE",x"FE",x"3B", -- 0x0108
		x"F4",x"EE",x"CD",x"54",x"83",x"08",x"44",x"55", -- 0x0110
		x"9A",x"82",x"21",x"55",x"24",x"A9",x"4B",x"55", -- 0x0118
		x"DF",x"AE",x"51",x"23",x"81",x"16",x"AF",x"F5", -- 0x0120
		x"E4",x"A2",x"50",x"B8",x"9C",x"9D",x"0F",x"6C", -- 0x0128
		x"FC",x"FE",x"7D",x"F5",x"B1",x"52",x"4C",x"ED", -- 0x0130
		x"8A",x"FA",x"31",x"75",x"66",x"EB",x"AB",x"D5", -- 0x0138
		x"FC",x"34",x"49",x"31",x"47",x"1E",x"3C",x"FA", -- 0x0140
		x"D4",x"AA",x"68",x"33",x"69",x"96",x"D4",x"2B", -- 0x0148
		x"F4",x"AA",x"E9",x"54",x"83",x"88",x"44",x"55", -- 0x0150
		x"9A",x"82",x"21",x"55",x"66",x"8B",x"EB",x"55", -- 0x0158
		x"FE",x"DC",x"DD",x"A9",x"90",x"EA",x"63",x"01", -- 0x0160
		x"88",x"F5",x"D3",x"C9",x"43",x"A0",x"98",x"FF", -- 0x0168
		x"F4",x"6E",x"25",x"33",x"BF",x"FF",x"FF",x"7D", -- 0x0170
		x"4B",x"A3",x"8D",x"17",x"C7",x"0D",x"C1",x"F3", -- 0x0178
		x"AA",x"54",x"95",x"EA",x"5A",x"35",x"95",x"9A", -- 0x0180
		x"CC",x"FA",x"7B",x"4D",x"63",x"99",x"AC",x"4E", -- 0x0188
		x"B4",x"AE",x"4D",x"55",x"A3",x"AA",x"44",x"55", -- 0x0190
		x"9A",x"8A",x"25",x"55",x"24",x"0B",x"AB",x"D5", -- 0x0198
		x"EF",x"47",x"13",x"11",x"C8",x"7E",x"7F",x"BB", -- 0x01A0
		x"DF",x"3E",x"7C",x"F3",x"E9",x"94",x"DA",x"2B", -- 0x01A8
		x"FC",x"7E",x"FD",x"D4",x"83",x"48",x"C4",x"D5", -- 0x01B0
		x"9A",x"82",x"21",x"55",x"62",x"A9",x"AB",x"55", -- 0x01B8
		x"3F",x"DF",x"6C",x"F3",x"FA",x"AD",x"BB",x"D3", -- 0x01C0
		x"DF",x"E5",x"F1",x"4C",x"F2",x"EA",x"77",x"BD", -- 0x01C8
		x"F7",x"AB",x"DB",x"65",x"52",x"05",x"AE",x"D9", -- 0x01D0
		x"E1",x"41",x"03",x"13",x"7A",x"FF",x"EB",x"D5", -- 0x01D8
		x"AA",x"34",x"FD",x"CE",x"C3",x"DC",x"5E",x"6E", -- 0x01E0
		x"AE",x"F8",x"6D",x"1E",x"4E",x"17",x"81",x"E3", -- 0x01E8
		x"B4",x"A2",x"4F",x"39",x"E0",x"EC",x"CF",x"86", -- 0x01F0
		x"4B",x"55",x"E2",x"FB",x"67",x"19",x"14",x"FF", -- 0x01F8
		x"AA",x"54",x"51",x"AB",x"2F",x"7F",x"DD",x"ED", -- 0x0200
		x"1B",x"B9",x"5C",x"5E",x"6C",x"96",x"AB",x"4F", -- 0x0208
		x"B4",x"BE",x"71",x"C5",x"FE",x"DF",x"D7",x"CD", -- 0x0210
		x"AE",x"7D",x"B7",x"BF",x"9B",x"06",x"A9",x"CF", -- 0x0218
		x"AA",x"54",x"55",x"AA",x"2A",x"C5",x"AD",x"2A", -- 0x0220
		x"D4",x"AA",x"6B",x"52",x"48",x"93",x"D3",x"2B", -- 0x0228
		x"B4",x"AE",x"4D",x"55",x"A3",x"AA",x"45",x"57", -- 0x0230
		x"9C",x"B2",x"45",x"6A",x"ED",x"DF",x"C9",x"9B", -- 0x0238
		x"AB",x"57",x"44",x"AF",x"2D",x"D1",x"B3",x"38", -- 0x0240
		x"DC",x"BC",x"79",x"53",x"37",x"BF",x"DC",x"3B", -- 0x0248
		x"09",x"13",x"D5",x"E1",x"E2",x"73",x"5D",x"AB", -- 0x0250
		x"7F",x"37",x"37",x"9B",x"6A",x"B5",x"5F",x"27", -- 0x0258
		x"B0",x"7A",x"7B",x"C1",x"C7",x"8A",x"E5",x"CC", -- 0x0260
		x"D7",x"87",x"49",x"4B",x"67",x"A2",x"D1",x"39", -- 0x0268
		x"5F",x"E7",x"AB",x"BF",x"DF",x"BD",x"17",x"6B", -- 0x0270
		x"FF",x"B7",x"37",x"9B",x"6A",x"75",x"DF",x"27", -- 0x0278
		x"B8",x"59",x"51",x"B8",x"18",x"DC",x"AC",x"2C", -- 0x0280
		x"D6",x"89",x"4B",x"13",x"25",x"82",x"D3",x"3B", -- 0x0288
		x"DF",x"E7",x"6B",x"27",x"FF",x"7D",x"57",x"2B", -- 0x0290
		x"47",x"03",x"17",x"9B",x"EA",x"95",x"1F",x"27", -- 0x0298
		x"AB",x"54",x"45",x"AA",x"2A",x"D5",x"AD",x"2A", -- 0x02A0
		x"D4",x"AA",x"49",x"12",x"65",x"96",x"DA",x"2B", -- 0x02A8
		x"D9",x"D3",x"B5",x"41",x"C2",x"A3",x"58",x"56", -- 0x02B0
		x"9B",x"AB",x"25",x"55",x"22",x"A9",x"AB",x"55", -- 0x02B8
		x"FF",x"5E",x"17",x"96",x"C8",x"77",x"1F",x"06", -- 0x02C0
		x"CE",x"E7",x"63",x"30",x"50",x"9C",x"8A",x"2B", -- 0x02C8
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"D7",x"EB", -- 0x02D0
		x"FF",x"77",x"77",x"DB",x"6A",x"55",x"5F",x"27", -- 0x02D8
		x"EE",x"47",x"17",x"11",x"DB",x"02",x"44",x"E1", -- 0x02E0
		x"F4",x"BB",x"57",x"3B",x"65",x"96",x"DA",x"2B", -- 0x02E8
		x"19",x"3E",x"2F",x"E5",x"43",x"E4",x"9C",x"FC", -- 0x02F0
		x"FB",x"CB",x"A5",x"55",x"36",x"D9",x"AB",x"55", -- 0x02F8
		x"AA",x"54",x"D1",x"F8",x"3B",x"EF",x"BD",x"78", -- 0x0300
		x"9D",x"74",x"EF",x"36",x"70",x"29",x"BF",x"EF", -- 0x0308
		x"B4",x"AA",x"4B",x"54",x"EB",x"1C",x"CD",x"EF", -- 0x0310
		x"67",x"FF",x"AE",x"CF",x"C7",x"69",x"34",x"FF", -- 0x0318
		x"AA",x"54",x"55",x"AA",x"2A",x"D5",x"AF",x"AF", -- 0x0320
		x"5F",x"9E",x"4F",x"27",x"72",x"3B",x"9F",x"CF", -- 0x0328
		x"B4",x"AE",x"4D",x"55",x"AB",x"FA",x"8D",x"E7", -- 0x0330
		x"F7",x"D7",x"E6",x"FB",x"A7",x"49",x"14",x"FF", -- 0x0338
		x"EE",x"47",x"15",x"56",x"E9",x"6C",x"65",x"C3", -- 0x0340
		x"E1",x"BF",x"5F",x"57",x"25",x"92",x"D6",x"2B", -- 0x0348
		x"97",x"0B",x"1B",x"85",x"E2",x"D9",x"CF",x"F1", -- 0x0350
		x"22",x"71",x"A8",x"54",x"67",x"A9",x"AB",x"55", -- 0x0358
		x"EF",x"52",x"19",x"83",x"85",x"C3",x"EF",x"3F", -- 0x0360
		x"DC",x"AA",x"68",x"53",x"6D",x"92",x"D6",x"2B", -- 0x0368
		x"E9",x"C6",x"EF",x"E3",x"65",x"20",x"5E",x"57", -- 0x0370
		x"9B",x"83",x"21",x"55",x"66",x"AB",x"AB",x"55", -- 0x0378
		x"53",x"96",x"AD",x"6A",x"AA",x"92",x"5E",x"2C", -- 0x0380
		x"56",x"57",x"AB",x"AB",x"AD",x"55",x"57",x"6B", -- 0x0388
		x"9F",x"27",x"2B",x"9F",x"97",x"2D",x"17",x"6B", -- 0x0390
		x"3B",x"17",x"35",x"9B",x"EA",x"35",x"1F",x"A7", -- 0x0398
		x"57",x"A8",x"B0",x"60",x"F8",x"6C",x"F4",x"EF", -- 0x03A0
		x"FF",x"7F",x"FD",x"FF",x"BF",x"7D",x"4B",x"D4", -- 0x03A8
		x"EB",x"59",x"36",x"1B",x"04",x"03",x"03",x"02", -- 0x03B0
		x"C5",x"F5",x"BA",x"FA",x"ED",x"B6",x"58",x"AA", -- 0x03B8
		x"55",x"2B",x"2E",x"1F",x"FD",x"2C",x"7C",x"DE", -- 0x03C0
		x"7E",x"7F",x"FF",x"BE",x"9F",x"77",x"2B",x"D4", -- 0x03C8
		x"4B",x"B5",x"AA",x"CA",x"F6",x"75",x"3F",x"3E", -- 0x03D0
		x"9D",x"1D",x"3A",x"FA",x"FD",x"D6",x"54",x"AA", -- 0x03D8
		x"B3",x"E9",x"DF",x"54",x"AE",x"AD",x"FF",x"7F", -- 0x03E0
		x"9F",x"DE",x"2F",x"AB",x"D3",x"55",x"BB",x"C9", -- 0x03E8
		x"F5",x"EB",x"3C",x"17",x"0D",x"0C",x"46",x"87", -- 0x03F0
		x"A5",x"C7",x"EE",x"F5",x"ED",x"EA",x"37",x"D9", -- 0x03F8
		x"F8",x"FE",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF", -- 0x0400
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0408
		x"7F",x"3F",x"3F",x"3F",x"8F",x"07",x"A3",x"D0", -- 0x0410
		x"E0",x"FA",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0418
		x"1F",x"8F",x"E7",x"E2",x"F9",x"FD",x"F8",x"FC", -- 0x0420
		x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0428
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"DE", -- 0x0430
		x"70",x"10",x"02",x"A3",x"CF",x"FF",x"FF",x"FF", -- 0x0438
		x"FF",x"FF",x"FF",x"3F",x"1F",x"07",x"82",x"43", -- 0x0440
		x"D0",x"E0",x"F8",x"FC",x"FF",x"FF",x"FF",x"FF", -- 0x0448
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC", -- 0x0450
		x"E4",x"00",x"04",x"93",x"5F",x"7F",x"FF",x"FF", -- 0x0458
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3E", -- 0x0460
		x"0F",x"01",x"40",x"E0",x"DA",x"FF",x"FF",x"FF", -- 0x0468
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EC", -- 0x0470
		x"F8",x"41",x"00",x"4B",x"0F",x"7F",x"FF",x"FF", -- 0x0478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0480
		x"FF",x"FF",x"FF",x"3F",x"16",x"42",x"C0",x"FF", -- 0x0488
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC", -- 0x0490
		x"F4",x"E1",x"84",x"0B",x"0F",x"3F",x"BF",x"FF", -- 0x0498
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04A0
		x"FF",x"FF",x"FF",x"FF",x"F9",x"C0",x"03",x"7F", -- 0x04A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC", -- 0x04B0
		x"F8",x"E0",x"C5",x"43",x"0F",x"3F",x"FF",x"FF", -- 0x04B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04C0
		x"FF",x"FF",x"FF",x"FE",x"F8",x"F0",x"F1",x"C2", -- 0x04C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC", -- 0x04D0
		x"F0",x"C0",x"82",x"13",x"1F",x"7F",x"FF",x"FF", -- 0x04D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x04E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EC", -- 0x04F0
		x"F0",x"E0",x"C5",x"83",x"0F",x"2F",x"1F",x"1F", -- 0x04F8
		x"FF",x"FF",x"FF",x"3F",x"0F",x"0B",x"84",x"20", -- 0x0500
		x"C0",x"F4",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0508
		x"FF",x"FF",x"FF",x"FC",x"F0",x"D0",x"42",x"04", -- 0x0510
		x"23",x"8F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0520
		x"FF",x"FF",x"FF",x"3F",x"0E",x"80",x"E0",x"FF", -- 0x0528
		x"FF",x"FF",x"FF",x"FC",x"F4",x"F0",x"E1",x"C2", -- 0x0530
		x"CB",x"87",x"8F",x"2F",x"3F",x"7F",x"BF",x"FF", -- 0x0538
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD", -- 0x0540
		x"FE",x"F8",x"E1",x"C5",x"8B",x"9F",x"3F",x"7F", -- 0x0548
		x"FF",x"FF",x"FF",x"FC",x"F8",x"F0",x"C2",x"80", -- 0x0550
		x"13",x"1F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0558
		x"1F",x"87",x"C3",x"F4",x"F8",x"FE",x"FE",x"FF", -- 0x0560
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0568
		x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"BF", -- 0x0570
		x"1F",x"9F",x"8F",x"CC",x"C0",x"E9",x"F3",x"FF", -- 0x0578
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0580
		x"FF",x"FF",x"FF",x"3F",x"0F",x"81",x"E8",x"FF", -- 0x0588
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0590
		x"FF",x"FF",x"FF",x"FC",x"E0",x"09",x"07",x"FF", -- 0x0598
		x"FF",x"FF",x"FE",x"FF",x"FE",x"FC",x"FD",x"FE", -- 0x05A0
		x"FC",x"FC",x"FD",x"FF",x"FE",x"FE",x"FF",x"FF", -- 0x05A8
		x"87",x"C7",x"4F",x"0F",x"1F",x"1F",x"1F",x"1F", -- 0x05B0
		x"BF",x"1F",x"3F",x"0F",x"0F",x"97",x"C7",x"03", -- 0x05B8
		x"F8",x"FC",x"F0",x"F4",x"F1",x"E1",x"F1",x"E3", -- 0x05C0
		x"E9",x"F1",x"E3",x"F8",x"F0",x"F4",x"F8",x"F8", -- 0x05C8
		x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F", -- 0x05D8
		x"CB",x"C7",x"8F",x"AF",x"8F",x"9F",x"9F",x"9F", -- 0x05E0
		x"9F",x"9F",x"9F",x"8F",x"CF",x"8F",x"E7",x"C7", -- 0x05E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F8
		x"FF",x"FF",x"FE",x"FE",x"FF",x"FE",x"FF",x"FF", -- 0x0600
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0608
		x"87",x"27",x"0F",x"8F",x"0F",x"1F",x"1F",x"4F", -- 0x0610
		x"87",x"A7",x"B3",x"E1",x"F9",x"F8",x"F8",x"FE", -- 0x0618
		x"FA",x"F8",x"F0",x"F8",x"C3",x"E9",x"F1",x"E0", -- 0x0620
		x"FA",x"FD",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0628
		x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0630
		x"FF",x"3F",x"07",x"C3",x"F1",x"F9",x"F8",x"FE", -- 0x0638
		x"C7",x"C7",x"CF",x"CF",x"C7",x"E7",x"E3",x"E0", -- 0x0640
		x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0650
		x"7F",x"0F",x"83",x"E3",x"F1",x"F8",x"F8",x"FE", -- 0x0658
		x"3F",x"9F",x"CF",x"CF",x"C7",x"E7",x"F7",x"E3", -- 0x0660
		x"EB",x"F1",x"F0",x"FA",x"FC",x"FF",x"FF",x"FF", -- 0x0668
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0670
		x"FF",x"FF",x"7F",x"3F",x"07",x"83",x"B8",x"FE", -- 0x0678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0680
		x"FF",x"FF",x"FF",x"FC",x"F8",x"F0",x"E1",x"C2", -- 0x0688
		x"FC",x"F9",x"F3",x"F3",x"F3",x"E7",x"E7",x"C3", -- 0x0690
		x"E7",x"CF",x"0F",x"1F",x"3F",x"7F",x"FF",x"FF", -- 0x0698
		x"C7",x"A7",x"CF",x"AF",x"9F",x"CF",x"E3",x"E0", -- 0x06A0
		x"F8",x"FA",x"FC",x"FE",x"FE",x"FF",x"FE",x"FF", -- 0x06A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06B0
		x"7F",x"3F",x"1F",x"9F",x"0F",x"8F",x"47",x"03", -- 0x06B8
		x"FA",x"F8",x"F4",x"F0",x"C9",x"E9",x"F1",x"F0", -- 0x06C0
		x"F4",x"F8",x"FD",x"FF",x"FE",x"FF",x"FE",x"FF", -- 0x06C8
		x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06D0
		x"7F",x"3F",x"3F",x"1F",x"8F",x"0F",x"4F",x"07", -- 0x06D8
		x"F8",x"FC",x"F0",x"F8",x"F1",x"E2",x"F1",x"C3", -- 0x06E0
		x"A3",x"8F",x"9F",x"9F",x"CF",x"8F",x"C7",x"C7", -- 0x06E8
		x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0700
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE", -- 0x0708
		x"FC",x"F9",x"F9",x"F9",x"F1",x"F1",x"F3",x"F3", -- 0x0710
		x"E3",x"E7",x"C7",x"87",x"1F",x"0F",x"5F",x"1F", -- 0x0718
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"9F", -- 0x0720
		x"8E",x"2E",x"0A",x"34",x"11",x"87",x"3A",x"0E", -- 0x0728
		x"48",x"C4",x"A2",x"C1",x"D3",x"E1",x"F7",x"66", -- 0x0730
		x"37",x"7B",x"F9",x"5B",x"62",x"BD",x"4B",x"A7", -- 0x0738
		x"2B",x"67",x"15",x"2A",x"26",x"09",x"1C",x"89", -- 0x0740
		x"83",x"C7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0748
		x"F7",x"AB",x"7B",x"B7",x"52",x"05",x"2F",x"1E", -- 0x0750
		x"8B",x"17",x"03",x"80",x"C1",x"E2",x"C4",x"08", -- 0x0758
		x"2E",x"DF",x"56",x"0B",x"D1",x"63",x"6F",x"3F", -- 0x0760
		x"DF",x"3F",x"1F",x"07",x"07",x"0B",x"23",x"12", -- 0x0768
		x"B9",x"2F",x"13",x"07",x"CF",x"FF",x"FF",x"FF", -- 0x0770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0788
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0790
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F8
		x"FF",x"CC",x"DA",x"A6",x"60",x"22",x"7F",x"FF", -- 0x0800
		x"7F",x"7F",x"7F",x"03",x"03",x"F3",x"F3",x"F3", -- 0x0808
		x"FF",x"29",x"D5",x"55",x"2D",x"09",x"19",x"C9", -- 0x0810
		x"C9",x"ED",x"C9",x"E5",x"D7",x"E9",x"C9",x"CD", -- 0x0818
		x"F3",x"F3",x"F3",x"F3",x"F3",x"F0",x"F1",x"FF", -- 0x0820
		x"FF",x"FF",x"FE",x"D9",x"74",x"38",x"04",x"4F", -- 0x0828
		x"F1",x"C3",x"ED",x"F9",x"A9",x"A5",x"19",x"39", -- 0x0830
		x"11",x"1D",x"95",x"3B",x"7F",x"2D",x"19",x"15", -- 0x0838
		x"FC",x"8A",x"80",x"20",x"40",x"28",x"0C",x"00", -- 0x0840
		x"00",x"18",x"22",x"18",x"08",x"03",x"07",x"E2", -- 0x0848
		x"09",x"8D",x"21",x"39",x"61",x"01",x"01",x"01", -- 0x0850
		x"19",x"15",x"29",x"0B",x"1F",x"15",x"2D",x"39", -- 0x0858
		x"CC",x"56",x"67",x"C2",x"80",x"D2",x"A4",x"9E", -- 0x0860
		x"F9",x"E3",x"31",x"18",x"08",x"00",x"FF",x"FF", -- 0x0868
		x"11",x"01",x"81",x"61",x"41",x"E1",x"B9",x"21", -- 0x0870
		x"99",x"99",x"21",x"61",x"21",x"01",x"FF",x"FF", -- 0x0878
		x"FF",x"EA",x"05",x"24",x"38",x"56",x"89",x"D4", -- 0x0880
		x"EE",x"A7",x"03",x"02",x"01",x"05",x"06",x"06", -- 0x0888
		x"FF",x"77",x"2F",x"33",x"5B",x"3D",x"D7",x"AB", -- 0x0890
		x"DB",x"55",x"77",x"FB",x"69",x"DB",x"E3",x"E7", -- 0x0898
		x"1E",x"0D",x"05",x"04",x"00",x"02",x"04",x"06", -- 0x08A0
		x"0F",x"07",x"07",x"01",x"43",x"40",x"69",x"B7", -- 0x08A8
		x"E3",x"63",x"35",x"2D",x"13",x"03",x"03",x"C5", -- 0x08B0
		x"43",x"51",x"33",x"DF",x"57",x"E7",x"E5",x"F1", -- 0x08B8
		x"DB",x"3E",x"37",x"04",x"00",x"C6",x"A9",x"54", -- 0x08C0
		x"6E",x"27",x"43",x"02",x"01",x"05",x"16",x"0E", -- 0x08C8
		x"5F",x"67",x"01",x"03",x"57",x"31",x"DB",x"CB", -- 0x08D0
		x"CD",x"77",x"63",x"D3",x"63",x"59",x"9B",x"E5", -- 0x08D8
		x"1F",x"05",x"01",x"4C",x"70",x"22",x"74",x"3A", -- 0x08E0
		x"0E",x"07",x"07",x"00",x"00",x"D3",x"FF",x"FF", -- 0x08E8
		x"ED",x"5F",x"1F",x"29",x"03",x"83",x"C1",x"D1", -- 0x08F0
		x"F3",x"DB",x"3F",x"11",x"03",x"17",x"FF",x"FF", -- 0x08F8
		x"FF",x"C2",x"C4",x"CF",x"C4",x"C9",x"CB",x"C7", -- 0x0900
		x"DB",x"C2",x"DA",x"8E",x"9E",x"C5",x"DF",x"C7", -- 0x0908
		x"FF",x"0C",x"1A",x"15",x"84",x"61",x"FF",x"FF", -- 0x0910
		x"7F",x"7E",x"7E",x"06",x"0E",x"FF",x"FF",x"FF", -- 0x0918
		x"9D",x"CF",x"D3",x"F9",x"8B",x"F9",x"9A",x"9B", -- 0x0920
		x"BF",x"8A",x"C6",x"DD",x"CC",x"C5",x"CE",x"CB", -- 0x0928
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x0930
		x"FF",x"FF",x"BF",x"67",x"97",x"03",x"05",x"87", -- 0x0938
		x"C7",x"C0",x"C0",x"C0",x"C0",x"D4",x"84",x"94", -- 0x0940
		x"88",x"9C",x"CB",x"CC",x"86",x"8B",x"C2",x"C1", -- 0x0948
		x"0B",x"47",x"80",x"40",x"D0",x"72",x"23",x"21", -- 0x0950
		x"4A",x"0C",x"BE",x"17",x"8F",x"C3",x"C2",x"80", -- 0x0958
		x"C7",x"C5",x"D2",x"D5",x"CB",x"C9",x"C5",x"C4", -- 0x0960
		x"C2",x"C1",x"CA",x"C1",x"C0",x"C0",x"FF",x"FF", -- 0x0968
		x"58",x"B9",x"1C",x"15",x"CF",x"A2",x"71",x"91", -- 0x0970
		x"0F",x"85",x"9B",x"02",x"00",x"00",x"C7",x"FF", -- 0x0978
		x"FF",x"F8",x"E7",x"C4",x"C0",x"E6",x"CB",x"F4", -- 0x0980
		x"CC",x"CF",x"C7",x"C2",x"E0",x"E0",x"E0",x"DC", -- 0x0988
		x"FF",x"04",x"0A",x"D8",x"4D",x"05",x"C5",x"AB", -- 0x0990
		x"DF",x"57",x"75",x"F0",x"D8",x"48",x"00",x"00", -- 0x0998
		x"E5",x"CE",x"CA",x"C7",x"E2",x"E0",x"F0",x"C2", -- 0x09A0
		x"E1",x"E2",x"C6",x"E0",x"C2",x"EC",x"E7",x"CF", -- 0x09A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x09B0
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09B8
		x"C7",x"E2",x"E0",x"C0",x"E0",x"E0",x"D6",x"C7", -- 0x09C0
		x"E4",x"E2",x"F2",x"D4",x"E2",x"E1",x"C7",x"E7", -- 0x09C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x09D0
		x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"00", -- 0x09D8
		x"E4",x"E0",x"CE",x"C5",x"E3",x"E0",x"C0",x"E0", -- 0x09E0
		x"E0",x"E0",x"C0",x"C0",x"E8",x"F3",x"FF",x"FF", -- 0x09E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04", -- 0x09F0
		x"0D",x"05",x"00",x"00",x"42",x"AE",x"FF",x"FF", -- 0x09F8
		x"FF",x"C0",x"DF",x"DF",x"DF",x"C0",x"CE",x"CE", -- 0x0A00
		x"CE",x"CE",x"C1",x"C1",x"DD",x"DD",x"DD",x"DF", -- 0x0A08
		x"FF",x"02",x"86",x"8C",x"99",x"11",x"33",x"67", -- 0x0A10
		x"C7",x"8F",x"9E",x"1E",x"3C",x"3C",x"39",x"31", -- 0x0A18
		x"C2",x"C6",x"C4",x"C4",x"C4",x"C4",x"CC",x"C9", -- 0x0A20
		x"C9",x"D9",x"D1",x"D1",x"D3",x"DF",x"DF",x"F0", -- 0x0A28
		x"70",x"60",x"60",x"E7",x"E7",x"C7",x"C7",x"C7", -- 0x0A30
		x"C1",x"CD",x"CD",x"8D",x"81",x"FF",x"FF",x"21", -- 0x0A38
		x"E3",x"E7",x"E6",x"E6",x"E6",x"C6",x"CE",x"CC", -- 0x0A40
		x"CC",x"DC",x"DC",x"9C",x"39",x"39",x"39",x"73", -- 0x0A48
		x"2F",x"2F",x"6F",x"4F",x"41",x"4F",x"4F",x"CF", -- 0x0A50
		x"8F",x"8F",x"8F",x"8F",x"8F",x"0F",x"01",x"1D", -- 0x0A58
		x"72",x"72",x"F7",x"E7",x"E4",x"C4",x"8F",x"9B", -- 0x0A60
		x"33",x"7B",x"58",x"DF",x"DF",x"C0",x"FF",x"FF", -- 0x0A68
		x"1D",x"01",x"FF",x"FF",x"1F",x"1F",x"9F",x"9F", -- 0x0A70
		x"9F",x"9F",x"1F",x"DF",x"C1",x"01",x"FF",x"FF", -- 0x0A78
		x"FF",x"DE",x"DE",x"DF",x"C3",x"FE",x"FF",x"CF", -- 0x0A80
		x"CF",x"CF",x"C0",x"C1",x"DD",x"DD",x"DD",x"C0", -- 0x0A88
		x"FF",x"07",x"3F",x"F9",x"DF",x"1F",x"9F",x"9F", -- 0x0A90
		x"9F",x"81",x"0F",x"CF",x"CF",x"CF",x"C1",x"01", -- 0x0A98
		x"DE",x"FE",x"E0",x"CE",x"CE",x"CE",x"CE",x"C0", -- 0x0AA0
		x"C0",x"FF",x"FF",x"CF",x"CF",x"CE",x"CE",x"C0", -- 0x0AA8
		x"F7",x"F7",x"F7",x"F7",x"01",x"DF",x"FF",x"FF", -- 0x0AB0
		x"21",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"0F", -- 0x0AB8
		x"C0",x"DC",x"DE",x"DE",x"DE",x"DE",x"C0",x"FC", -- 0x0AC0
		x"FE",x"C7",x"C0",x"DE",x"DE",x"DF",x"DF",x"DF", -- 0x0AC8
		x"01",x"01",x"01",x"07",x"07",x"07",x"E7",x"E7", -- 0x0AD0
		x"07",x"F1",x"E1",x"01",x"DF",x"DF",x"DF",x"DF", -- 0x0AD8
		x"DF",x"C1",x"C0",x"CF",x"CF",x"CF",x"CF",x"CF", -- 0x0AE0
		x"C0",x"C0",x"C7",x"C7",x"C7",x"C0",x"FF",x"FF", -- 0x0AE8
		x"C1",x"3D",x"3D",x"BD",x"81",x"9F",x"BF",x"A1", -- 0x0AF0
		x"1F",x"1F",x"9F",x"9F",x"9F",x"01",x"FF",x"FF", -- 0x0AF8
		x"FF",x"F7",x"BF",x"B8",x"B7",x"BF",x"BF",x"88", -- 0x0B00
		x"FF",x"FF",x"FF",x"DC",x"DC",x"DC",x"DC",x"DC", -- 0x0B08
		x"FF",x"3F",x"3F",x"3F",x"3F",x"3F",x"01",x"01", -- 0x0B10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B18
		x"C0",x"CE",x"CE",x"CF",x"CF",x"CF",x"C1",x"C1", -- 0x0B20
		x"CF",x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"CF", -- 0x0B28
		x"01",x"1F",x"DF",x"DF",x"C1",x"DF",x"FF",x"21", -- 0x0B30
		x"3F",x"3F",x"3F",x"3F",x"3F",x"01",x"01",x"BF", -- 0x0B38
		x"CF",x"CF",x"CC",x"CC",x"CD",x"CF",x"CF",x"CE", -- 0x0B40
		x"C0",x"C7",x"FF",x"FC",x"CF",x"CF",x"CF",x"C0", -- 0x0B48
		x"BF",x"BF",x"3F",x"3F",x"BF",x"BF",x"81",x"07", -- 0x0B50
		x"FF",x"F1",x"8F",x"6F",x"EF",x"EF",x"EF",x"8F", -- 0x0B58
		x"C0",x"DF",x"DF",x"DF",x"DF",x"C0",x"CF",x"CF", -- 0x0B60
		x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF", -- 0x0B68
		x"61",x"6F",x"7F",x"7F",x"71",x"1F",x"9F",x"9F", -- 0x0B70
		x"9F",x"9F",x"9F",x"9F",x"01",x"01",x"FF",x"FF", -- 0x0B78
		x"FF",x"C0",x"DE",x"DE",x"DE",x"DE",x"DE",x"DE", -- 0x0B80
		x"C0",x"DF",x"DF",x"DF",x"DF",x"C0",x"FF",x"FF", -- 0x0B88
		x"FF",x"1B",x"61",x"75",x"39",x"1F",x"17",x"05", -- 0x0B90
		x"19",x"15",x"0D",x"27",x"3F",x"0D",x"27",x"FF", -- 0x0B98
		x"FF",x"DB",x"DF",x"DF",x"DF",x"DF",x"DF",x"C4", -- 0x0BA0
		x"DE",x"DE",x"DF",x"DF",x"C0",x"DE",x"DE",x"DE", -- 0x0BA8
		x"FF",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"01", -- 0x0BB0
		x"01",x"C1",x"E1",x"21",x"E1",x"E1",x"E1",x"E1", -- 0x0BB8
		x"DE",x"C0",x"CF",x"CF",x"CF",x"CF",x"CF",x"C0", -- 0x0BC0
		x"C0",x"CF",x"FF",x"FE",x"CE",x"CE",x"CE",x"C0", -- 0x0BC8
		x"E1",x"07",x"7F",x"7F",x"7F",x"7F",x"79",x"01", -- 0x0BD0
		x"1F",x"FF",x"FF",x"0F",x"EF",x"EF",x"E1",x"E1", -- 0x0BD8
		x"C0",x"DE",x"FE",x"FE",x"FF",x"E1",x"CF",x"CF", -- 0x0BE0
		x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF", -- 0x0BE8
		x"EF",x"0F",x"0F",x"EF",x"EF",x"01",x"81",x"9F", -- 0x0BF0
		x"9F",x"9F",x"9F",x"9F",x"01",x"01",x"FF",x"FF", -- 0x0BF8
		x"FF",x"CF",x"DB",x"DB",x"F3",x"F0",x"7E",x"5F", -- 0x0C00
		x"DF",x"DF",x"9E",x"81",x"BF",x"BF",x"80",x"9B", -- 0x0C08
		x"FF",x"CF",x"CF",x"CF",x"CF",x"01",x"C1",x"DF", -- 0x0C10
		x"DF",x"1F",x"C1",x"DF",x"DF",x"01",x"7D",x"7D", -- 0x0C18
		x"9B",x"80",x"FF",x"FF",x"B3",x"B3",x"B3",x"B3", -- 0x0C20
		x"83",x"B3",x"B0",x"B0",x"B0",x"80",x"FF",x"FF", -- 0x0C28
		x"7D",x"7D",x"07",x"FF",x"BF",x"BF",x"BF",x"BF", -- 0x0C30
		x"87",x"87",x"67",x"67",x"61",x"61",x"3F",x"FF", -- 0x0C38
		x"FF",x"00",x"FE",x"FE",x"FE",x"00",x"1E",x"FE", -- 0x0C40
		x"FE",x"FE",x"E1",x"0F",x"7E",x"F0",x"8F",x"0F", -- 0x0C48
		x"FF",x"01",x"07",x"0F",x"0F",x"79",x"79",x"79", -- 0x0C50
		x"07",x"1F",x"F9",x"C1",x"6D",x"7D",x"7D",x"71", -- 0x0C58
		x"EF",x"EF",x"E0",x"FD",x"1F",x"02",x"63",x"63", -- 0x0C60
		x"63",x"03",x"E3",x"E3",x"E0",x"00",x"FF",x"FF", -- 0x0C68
		x"1F",x"1F",x"1F",x"DF",x"DF",x"01",x"C7",x"C7", -- 0x0C70
		x"C1",x"CF",x"DF",x"DF",x"1F",x"11",x"FF",x"FF", -- 0x0C78
		x"FF",x"09",x"E3",x"E3",x"E3",x"E3",x"06",x"0F", -- 0x0C80
		x"FF",x"FD",x"8D",x"9D",x"99",x"18",x"FF",x"FF", -- 0x0C88
		x"FF",x"F7",x"7F",x"7F",x"7F",x"09",x"EF",x"FF", -- 0x0C90
		x"11",x"BF",x"BF",x"BF",x"BF",x"01",x"FF",x"FF", -- 0x0C98
		x"FF",x"F7",x"FF",x"F8",x"F7",x"07",x"07",x"E7", -- 0x0CA0
		x"E7",x"E0",x"E0",x"E7",x"0F",x"08",x"FF",x"FF", -- 0x0CA8
		x"FF",x"3F",x"3F",x"3F",x"BF",x"81",x"81",x"A1", -- 0x0CB0
		x"A1",x"21",x"21",x"A1",x"81",x"01",x"FF",x"FF", -- 0x0CB8
		x"FF",x"00",x"CE",x"DE",x"DE",x"DE",x"D0",x"C0", -- 0x0CC0
		x"20",x"1B",x"1F",x"33",x"17",x"03",x"84",x"F0", -- 0x0CC8
		x"FF",x"19",x"3D",x"5F",x"3F",x"2D",x"25",x"1F", -- 0x0CD0
		x"4F",x"1F",x"8B",x"C1",x"C1",x"41",x"7F",x"FF", -- 0x0CD8
		x"FF",x"0F",x"EF",x"EF",x"EF",x"E0",x"EE",x"0E", -- 0x0CE0
		x"0E",x"0E",x"01",x"1F",x"1F",x"01",x"FF",x"FF", -- 0x0CE8
		x"FF",x"BF",x"BF",x"BF",x"BF",x"01",x"EF",x"FF", -- 0x0CF0
		x"11",x"DF",x"DF",x"DF",x"DF",x"01",x"FF",x"FF", -- 0x0CF8
		x"FF",x"CE",x"CE",x"CE",x"CF",x"CF",x"C0",x"C0", -- 0x0D00
		x"FF",x"FF",x"DE",x"DE",x"DF",x"DF",x"DF",x"C1", -- 0x0D08
		x"FF",x"0F",x"0F",x"0F",x"FF",x"FF",x"00",x"00", -- 0x0D10
		x"FF",x"FF",x"07",x"F7",x"F7",x"F7",x"F7",x"07", -- 0x0D18
		x"DD",x"DD",x"DD",x"DD",x"DC",x"C0",x"DC",x"DC", -- 0x0D20
		x"DC",x"C0",x"DC",x"DC",x"DC",x"C0",x"FF",x"FF", -- 0x0D28
		x"E0",x"E0",x"E0",x"F0",x"10",x"F0",x"F0",x"F0", -- 0x0D30
		x"F0",x"EF",x"EF",x"E0",x"0E",x"0E",x"E3",x"FF", -- 0x0D38
		x"FF",x"DF",x"DF",x"DF",x"DF",x"C0",x"DE",x"DE", -- 0x0D40
		x"DF",x"DF",x"C0",x"DE",x"FE",x"FE",x"FE",x"E0", -- 0x0D48
		x"FF",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"F7", -- 0x0D50
		x"F7",x"07",x"F7",x"F0",x"F0",x"F3",x"1F",x"FC", -- 0x0D58
		x"C7",x"FD",x"F9",x"C1",x"C1",x"C0",x"E0",x"E1", -- 0x0D60
		x"E3",x"E2",x"E0",x"E1",x"E1",x"E1",x"FF",x"FF", -- 0x0D68
		x"FB",x"FB",x"FB",x"FB",x"F8",x"0B",x"0F",x"EF", -- 0x0D70
		x"EF",x"0C",x"FB",x"FB",x"FB",x"F8",x"1F",x"FF", -- 0x0D78
		x"FF",x"CF",x"CF",x"CF",x"CF",x"C0",x"DB",x"DF", -- 0x0D80
		x"DF",x"DF",x"DC",x"DD",x"DF",x"C2",x"FF",x"FF", -- 0x0D88
		x"FF",x"F0",x"E7",x"E7",x"E7",x"67",x"E0",x"E0", -- 0x0D90
		x"FF",x"FF",x"67",x"EF",x"EF",x"68",x"FF",x"FF", -- 0x0D98
		x"FF",x"DC",x"FD",x"E1",x"DD",x"DD",x"DD",x"DD", -- 0x0DA0
		x"C0",x"CE",x"DE",x"D0",x"DE",x"DE",x"C3",x"FF", -- 0x0DA8
		x"FF",x"10",x"F6",x"F6",x"F6",x"F6",x"F0",x"F3", -- 0x0DB0
		x"13",x"F3",x"F3",x"F3",x"F0",x"10",x"FF",x"FF", -- 0x0DB8
		x"FF",x"DF",x"FF",x"E0",x"DC",x"DC",x"C1",x"D9", -- 0x0DC0
		x"F9",x"F9",x"E1",x"D9",x"D8",x"C0",x"FF",x"FF", -- 0x0DC8
		x"FF",x"7C",x"7C",x"7D",x"7D",x"01",x"C1",x"C1", -- 0x0DD0
		x"DF",x"DE",x"DE",x"DE",x"00",x"00",x"FF",x"FF", -- 0x0DD8
		x"FF",x"D8",x"D8",x"DB",x"DF",x"DF",x"C7",x"DF", -- 0x0DE0
		x"FC",x"E7",x"C7",x"C7",x"C0",x"C0",x"FF",x"FF", -- 0x0DE8
		x"FF",x"CC",x"7D",x"FF",x"B3",x"B3",x"9B",x"9A", -- 0x0DF0
		x"0C",x"FC",x"F6",x"F6",x"02",x"02",x"FF",x"FF", -- 0x0DF8
		x"FF",x"C1",x"D9",x"D9",x"D8",x"D8",x"DB",x"C3", -- 0x0E00
		x"F9",x"FF",x"CD",x"DD",x"DD",x"7D",x"30",x"18", -- 0x0E08
		x"FF",x"F7",x"FF",x"FF",x"0F",x"09",x"7D",x"7D", -- 0x0E10
		x"07",x"FF",x"F1",x"F7",x"F7",x"F7",x"07",x"07", -- 0x0E18
		x"0C",x"06",x"1E",x"15",x"18",x"0A",x"04",x"0C", -- 0x0E20
		x"00",x"00",x"01",x"01",x"00",x"00",x"FE",x"FF", -- 0x0E28
		x"F1",x"F7",x"07",x"87",x"C7",x"61",x"31",x"99", -- 0x0E30
		x"CD",x"D7",x"E3",x"71",x"AD",x"49",x"2F",x"FF", -- 0x0E38
		x"FF",x"03",x"3F",x"3F",x"3F",x"3F",x"3F",x"03", -- 0x0E40
		x"03",x"FF",x"FF",x"1F",x"9F",x"9F",x"9F",x"1F", -- 0x0E48
		x"FF",x"7D",x"7D",x"7D",x"7D",x"01",x"DF",x"DF", -- 0x0E50
		x"DF",x"DF",x"1F",x"01",x"6F",x"FF",x"FD",x"7D", -- 0x0E58
		x"9F",x"83",x"83",x"0F",x"EF",x"EF",x"EF",x"E2", -- 0x0E60
		x"02",x"7E",x"7E",x"7E",x"7E",x"03",x"FF",x"FF", -- 0x0E68
		x"7D",x"01",x"DF",x"DF",x"DF",x"1F",x"C1",x"DD", -- 0x0E70
		x"DD",x"DD",x"DD",x"DD",x"1D",x"01",x"FF",x"FF", -- 0x0E78
		x"FF",x"D9",x"D9",x"D9",x"D9",x"D9",x"C1",x"C0", -- 0x0E80
		x"CF",x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"DC", -- 0x0E88
		x"FF",x"FF",x"FF",x"87",x"87",x"87",x"87",x"01", -- 0x0E90
		x"01",x"3D",x"3D",x"3D",x"01",x"01",x"EF",x"EF", -- 0x0E98
		x"FC",x"FC",x"FC",x"E0",x"C0",x"DC",x"FC",x"DC", -- 0x0EA0
		x"DC",x"DF",x"DF",x"DF",x"C0",x"C0",x"FF",x"FF", -- 0x0EA8
		x"EF",x"EF",x"E1",x"ED",x"FD",x"1D",x"11",x"01", -- 0x0EB0
		x"1F",x"DF",x"DF",x"DF",x"01",x"01",x"FF",x"FF", -- 0x0EB8
		x"FF",x"DF",x"DF",x"DF",x"C0",x"DC",x"DD",x"DF", -- 0x0EC0
		x"DF",x"C2",x"C7",x"C7",x"C7",x"C7",x"C0",x"FF", -- 0x0EC8
		x"FF",x"7F",x"7F",x"7F",x"07",x"07",x"F7",x"F7", -- 0x0ED0
		x"F1",x"1D",x"9D",x"9D",x"9D",x"9D",x"01",x"8F", -- 0x0ED8
		x"FF",x"F1",x"B1",x"B1",x"B1",x"B1",x"B0",x"80", -- 0x0EE0
		x"DE",x"DE",x"C0",x"DE",x"FE",x"E0",x"FF",x"FF", -- 0x0EE8
		x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"09",x"01", -- 0x0EF0
		x"DF",x"DF",x"DF",x"DF",x"DF",x"01",x"FF",x"FF", -- 0x0EF8
		x"FF",x"DE",x"DF",x"C1",x"DF",x"DE",x"DE",x"DE", -- 0x0F00
		x"DE",x"C0",x"FF",x"FF",x"C0",x"CF",x"DF",x"DF", -- 0x0F08
		x"FF",x"EF",x"EF",x"EF",x"00",x"3F",x"3F",x"3F", -- 0x0F10
		x"00",x"00",x"FF",x"FF",x"1E",x"9F",x"9F",x"87", -- 0x0F18
		x"D0",x"C0",x"CE",x"CE",x"CE",x"CE",x"CE",x"CF", -- 0x0F20
		x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF", -- 0x0F28
		x"37",x"37",x"F7",x"F7",x"F0",x"07",x"FF",x"FF", -- 0x0F30
		x"0F",x"FF",x"F8",x"F7",x"07",x"00",x"FF",x"FF", -- 0x0F38
		x"FF",x"CA",x"C9",x"E4",x"9E",x"8B",x"86",x"C0", -- 0x0F40
		x"C1",x"FF",x"FF",x"DE",x"DE",x"DE",x"DE",x"C0", -- 0x0F48
		x"FF",x"4F",x"4F",x"CF",x"CF",x"40",x"5C",x"DC", -- 0x0F50
		x"C0",x"FF",x"FF",x"00",x"F7",x"F7",x"F7",x"F0", -- 0x0F58
		x"DE",x"DE",x"DE",x"DE",x"C0",x"CF",x"CF",x"CF", -- 0x0F60
		x"CF",x"C0",x"C0",x"CE",x"DE",x"D0",x"FF",x"FF", -- 0x0F68
		x"F3",x"F7",x"07",x"3C",x"3B",x"BB",x"BB",x"83", -- 0x0F70
		x"80",x"03",x"83",x"83",x"83",x"80",x"FF",x"FF", -- 0x0F78
		x"FF",x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"DC", -- 0x0F80
		x"DC",x"DC",x"C3",x"DB",x"DB",x"DB",x"D8",x"C3", -- 0x0F88
		x"FF",x"DF",x"FF",x"FF",x"FF",x"21",x"7D",x"7D", -- 0x0F90
		x"7D",x"01",x"F7",x"F7",x"F7",x"F7",x"07",x"81", -- 0x0F98
		x"DF",x"FF",x"E4",x"CF",x"CF",x"CF",x"CF",x"C0", -- 0x0FA0
		x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"FF",x"FF", -- 0x0FA8
		x"81",x"C1",x"41",x"C1",x"C1",x"9F",x"9F",x"1F", -- 0x0FB0
		x"DF",x"DF",x"C1",x"DF",x"3F",x"21",x"FF",x"FF", -- 0x0FB8
		x"FF",x"CC",x"CC",x"CF",x"CF",x"CC",x"C0",x"C0", -- 0x0FC0
		x"FF",x"FF",x"DC",x"FC",x"FC",x"E0",x"DC",x"DC", -- 0x0FC8
		x"FF",x"67",x"67",x"E7",x"E7",x"67",x"01",x"01", -- 0x0FD0
		x"FF",x"FF",x"7F",x"7F",x"7F",x"7F",x"01",x"01", -- 0x0FD8
		x"DD",x"C1",x"F1",x"F9",x"DC",x"CE",x"DF",x"FB", -- 0x0FE0
		x"F9",x"FB",x"FB",x"E3",x"C3",x"C0",x"FF",x"FF", -- 0x0FE8
		x"EF",x"EF",x"EF",x"E1",x"1F",x"1F",x"1F",x"9F", -- 0x0FF0
		x"C1",x"E7",x"FF",x"B9",x"9D",x"0F",x"FF",x"FF", -- 0x0FF8
		x"FF",x"C0",x"DE",x"DE",x"DE",x"DE",x"DE",x"C0", -- 0x1000
		x"C0",x"FF",x"FF",x"C1",x"C3",x"C3",x"C2",x"FF", -- 0x1008
		x"FF",x"81",x"81",x"81",x"BD",x"BD",x"81",x"9F", -- 0x1010
		x"90",x"90",x"96",x"FE",x"FE",x"FE",x"38",x"E0", -- 0x1018
		x"FF",x"C3",x"DF",x"DF",x"DF",x"C3",x"FF",x"FF", -- 0x1020
		x"C0",x"C0",x"CF",x"CF",x"CF",x"CF",x"C0",x"C0", -- 0x1028
		x"FF",x"01",x"19",x"19",x"19",x"19",x"01",x"9F", -- 0x1030
		x"F1",x"61",x"27",x"2F",x"2F",x"2F",x"29",x"3F", -- 0x1038
		x"FE",x"C3",x"DE",x"DE",x"DE",x"C0",x"FF",x"FF", -- 0x1040
		x"C1",x"DD",x"DD",x"DD",x"DD",x"C1",x"C1",x"FF", -- 0x1048
		x"0E",x"8E",x"8E",x"80",x"84",x"84",x"84",x"FF", -- 0x1050
		x"FF",x"81",x"BD",x"BD",x"BD",x"BD",x"87",x"80", -- 0x1058
		x"FF",x"C0",x"DF",x"DF",x"DF",x"DF",x"C0",x"C0", -- 0x1060
		x"DF",x"DF",x"DE",x"DE",x"DE",x"C6",x"FF",x"FF", -- 0x1068
		x"FF",x"C1",x"CD",x"CD",x"CD",x"CD",x"C1",x"C1", -- 0x1070
		x"C1",x"C3",x"02",x"06",x"0C",x"18",x"F8",x"FC", -- 0x1078
		x"3F",x"23",x"23",x"23",x"33",x"19",x"11",x"11", -- 0x1080
		x"71",x"F1",x"FD",x"EF",x"8F",x"8F",x"81",x"FF", -- 0x1088
		x"FF",x"03",x"7F",x"7E",x"7C",x"0C",x"18",x"18", -- 0x1090
		x"F8",x"F8",x"3C",x"3C",x"3C",x"00",x"08",x"F8", -- 0x1098
		x"FF",x"DB",x"FB",x"FB",x"FB",x"E3",x"FF",x"7F", -- 0x10A0
		x"60",x"6F",x"4F",x"4F",x"4F",x"41",x"41",x"7F", -- 0x10A8
		x"FF",x"01",x"67",x"7F",x"7F",x"7F",x"01",x"FF", -- 0x10B0
		x"40",x"40",x"FF",x"FF",x"79",x"F9",x"F9",x"8F", -- 0x10B8
		x"FF",x"84",x"B4",x"B6",x"B2",x"B3",x"82",x"FE", -- 0x10C0
		x"42",x"4E",x"4E",x"4E",x"4E",x"42",x"7F",x"FF", -- 0x10C8
		x"FC",x"E4",x"E4",x"E4",x"04",x"FC",x"00",x"00", -- 0x10D0
		x"1F",x"FD",x"FD",x"FD",x"FD",x"01",x"FF",x"FF", -- 0x10D8
		x"7F",x"40",x"5C",x"7C",x"7C",x"7C",x"60",x"FF", -- 0x10E0
		x"FF",x"81",x"BD",x"BD",x"BD",x"81",x"FF",x"FF", -- 0x10E8
		x"FC",x"BC",x"BC",x"BC",x"86",x"82",x"82",x"FE", -- 0x10F0
		x"03",x"01",x"39",x"39",x"39",x"01",x"FF",x"FF", -- 0x10F8
		x"3F",x"2F",x"2F",x"20",x"3F",x"FF",x"F8",x"79", -- 0x1100
		x"7B",x"7B",x"7A",x"02",x"82",x"82",x"FF",x"FF", -- 0x1108
		x"FF",x"07",x"0D",x"19",x"FF",x"EF",x"CF",x"81", -- 0x1110
		x"FF",x"FF",x"01",x"7D",x"7D",x"7D",x"07",x"FF", -- 0x1118
		x"03",x"FE",x"FE",x"83",x"83",x"83",x"80",x"87", -- 0x1120
		x"87",x"FE",x"FE",x"86",x"F6",x"F6",x"F7",x"9F", -- 0x1128
		x"FF",x"31",x"37",x"F7",x"F7",x"F7",x"37",x"F1", -- 0x1130
		x"F1",x"3D",x"3D",x"3D",x"3D",x"01",x"FF",x"FF", -- 0x1138
		x"1F",x"38",x"38",x"BF",x"BF",x"BB",x"82",x"82", -- 0x1140
		x"82",x"82",x"82",x"BA",x"FA",x"C2",x"FE",x"FE", -- 0x1148
		x"FF",x"7B",x"7B",x"7B",x"03",x"E3",x"7F",x"7F", -- 0x1150
		x"63",x"6F",x"6F",x"6F",x"6F",x"63",x"7F",x"7F", -- 0x1158
		x"FC",x"84",x"B5",x"B7",x"B7",x"B6",x"B6",x"86", -- 0x1160
		x"FF",x"FF",x"82",x"9E",x"9E",x"9E",x"82",x"FE", -- 0x1168
		x"7F",x"C3",x"FB",x"BB",x"3B",x"3B",x"3B",x"03", -- 0x1170
		x"FF",x"FF",x"1F",x"1F",x"03",x"1B",x"1F",x"0F", -- 0x1178
		x"00",x"FF",x"FF",x"2E",x"2E",x"2E",x"2E",x"2E", -- 0x1180
		x"20",x"20",x"20",x"3E",x"3E",x"02",x"02",x"02", -- 0x1188
		x"00",x"E0",x"E0",x"24",x"20",x"20",x"20",x"20", -- 0x1190
		x"20",x"F8",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x1198
		x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"00", -- 0x11A0
		x"03",x"07",x"07",x"04",x"00",x"00",x"00",x"00", -- 0x11A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x11B0
		x"D0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00", -- 0x11B8
		x"10",x"10",x"10",x"10",x"17",x"17",x"17",x"17", -- 0x11C0
		x"10",x"FF",x"FF",x"02",x"12",x"02",x"02",x"02", -- 0x11C8
		x"00",x"00",x"1E",x"1E",x"C3",x"80",x"80",x"80", -- 0x11D0
		x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x11D8
		x"02",x"02",x"3E",x"3E",x"3E",x"02",x"FF",x"FF", -- 0x11E0
		x"20",x"38",x"38",x"38",x"38",x"38",x"20",x"3F", -- 0x11E8
		x"00",x"00",x"00",x"06",x"06",x"06",x"F6",x"F0", -- 0x11F0
		x"FF",x"FF",x"E0",x"E0",x"00",x"88",x"80",x"80", -- 0x11F8
		x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"FF", -- 0x1200
		x"03",x"21",x"00",x"01",x"C5",x"CA",x"C7",x"C7", -- 0x1208
		x"00",x"60",x"24",x"52",x"1A",x"3E",x"14",x"00", -- 0x1210
		x"80",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"70", -- 0x1218
		x"C2",x"C8",x"CD",x"C2",x"C6",x"C3",x"C1",x"C7", -- 0x1220
		x"CF",x"C3",x"C6",x"C2",x"C2",x"C0",x"3C",x"70", -- 0x1228
		x"70",x"70",x"F0",x"F0",x"00",x"00",x"00",x"F8", -- 0x1230
		x"78",x"78",x"78",x"78",x"78",x"78",x"00",x"00", -- 0x1238
		x"58",x"3F",x"F7",x"A7",x"00",x"40",x"C0",x"00", -- 0x1240
		x"38",x"38",x"38",x"38",x"18",x"F8",x"F8",x"F8", -- 0x1248
		x"00",x"F8",x"F8",x"F8",x"38",x"38",x"38",x"38", -- 0x1250
		x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"00", -- 0x1258
		x"00",x"00",x"00",x"00",x"FE",x"FE",x"FE",x"81", -- 0x1260
		x"C7",x"65",x"E3",x"00",x"80",x"00",x"00",x"00", -- 0x1268
		x"00",x"18",x"38",x"1C",x"1C",x"34",x"0E",x"1E", -- 0x1270
		x"0E",x"9C",x"14",x"14",x"00",x"00",x"00",x"00", -- 0x1278
		x"00",x"C0",x"60",x"00",x"00",x"FF",x"FF",x"DF", -- 0x1280
		x"C0",x"C3",x"C1",x"C3",x"C3",x"C1",x"00",x"00", -- 0x1288
		x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF", -- 0x1290
		x"00",x"83",x"E7",x"C7",x"E9",x"77",x"EE",x"5E", -- 0x1298
		x"00",x"F8",x"F8",x"D8",x"C0",x"C3",x"C7",x"C1", -- 0x12A0
		x"CA",x"0C",x"1C",x"04",x"00",x"00",x"00",x"FF", -- 0x12A8
		x"1C",x"0C",x"50",x"68",x"B0",x"7C",x"FC",x"DC", -- 0x12B0
		x"58",x"E8",x"D0",x"20",x"2E",x"1B",x"07",x"83", -- 0x12B8
		x"FF",x"DF",x"C0",x"C0",x"C6",x"C2",x"C3",x"C0", -- 0x12C0
		x"C0",x"C1",x"C1",x"C0",x"00",x"31",x"5B",x"7C", -- 0x12C8
		x"85",x"9D",x"19",x"0C",x"3E",x"1E",x"1E",x"0C", -- 0x12D0
		x"BC",x"98",x"F8",x"EA",x"E7",x"56",x"9A",x"91", -- 0x12D8
		x"B7",x"2F",x"07",x"0A",x"00",x"00",x"01",x"FF", -- 0x12E0
		x"FF",x"DE",x"F6",x"2F",x"03",x"06",x"00",x"00", -- 0x12E8
		x"8B",x"08",x"00",x"00",x"07",x"3F",x"FF",x"FE", -- 0x12F0
		x"CF",x"07",x"07",x"2E",x"14",x"00",x"00",x"00", -- 0x12F8
		x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"FE", -- 0x1300
		x"00",x"00",x"9C",x"DE",x"EE",x"7E",x"FA",x"54", -- 0x1308
		x"00",x"00",x"00",x"00",x"80",x"FF",x"FF",x"FF", -- 0x1310
		x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"01", -- 0x1318
		x"38",x"00",x"1F",x"1F",x"80",x"80",x"80",x"80", -- 0x1320
		x"80",x"80",x"00",x"00",x"00",x"00",x"10",x"10", -- 0x1328
		x"01",x"01",x"11",x"11",x"11",x"11",x"19",x"19", -- 0x1330
		x"19",x"19",x"19",x"19",x"19",x"01",x"10",x"10", -- 0x1338
		x"1F",x"80",x"80",x"83",x"05",x"0B",x"02",x"01", -- 0x1340
		x"E0",x"EF",x"EF",x"EF",x"00",x"9C",x"D7",x"CF", -- 0x1348
		x"F1",x"03",x"02",x"81",x"F0",x"B3",x"83",x"81", -- 0x1350
		x"80",x"C0",x"E0",x"F0",x"F8",x"7F",x"3F",x"1F", -- 0x1358
		x"0E",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00", -- 0x1360
		x"9C",x"BA",x"DF",x"17",x"09",x"04",x"00",x"00", -- 0x1368
		x"00",x"00",x"00",x"00",x"FF",x"F7",x"EB",x"07", -- 0x1370
		x"4F",x"EB",x"F4",x"5B",x"20",x"01",x"00",x"00", -- 0x1378
		x"00",x"06",x"0F",x"17",x"0E",x"0B",x"17",x"0A", -- 0x1380
		x"00",x"06",x"07",x"07",x"02",x"01",x"06",x"0C", -- 0x1388
		x"00",x"00",x"53",x"BF",x"B6",x"5B",x"39",x"09", -- 0x1390
		x"01",x"01",x"00",x"FF",x"FF",x"F7",x"70",x"70", -- 0x1398
		x"06",x"06",x"03",x"00",x"00",x"00",x"00",x"1F", -- 0x13A0
		x"1F",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x13A8
		x"70",x"7F",x"7F",x"3E",x"01",x"01",x"01",x"E1", -- 0x13B0
		x"E1",x"E0",x"18",x"0C",x"5C",x"3E",x"2E",x"5F", -- 0x13B8
		x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x13C0
		x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E",x"1E", -- 0x13C8
		x"15",x"2D",x"3D",x"19",x"11",x"01",x"01",x"01", -- 0x13D0
		x"00",x"20",x"3F",x"3F",x"38",x"38",x"38",x"38", -- 0x13D8
		x"07",x"07",x"03",x"05",x"0B",x"07",x"06",x"09", -- 0x13E0
		x"0A",x"01",x"05",x"00",x"00",x"00",x"00",x"00", -- 0x13E8
		x"B8",x"38",x"B8",x"B8",x"F8",x"F8",x"F8",x"BF", -- 0x13F0
		x"BF",x"BE",x"78",x"2F",x"15",x"02",x"00",x"00", -- 0x13F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00", -- 0x1400
		x"BE",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1408
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F", -- 0x1410
		x"C0",x"7B",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1418
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1420
		x"FF",x"3F",x"C0",x"3E",x"00",x"00",x"00",x"00", -- 0x1428
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1430
		x"FF",x"FF",x"3F",x"80",x"7B",x"00",x"00",x"00", -- 0x1438
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1440
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1448
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1450
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1458
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1460
		x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"00", -- 0x1468
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1470
		x"00",x"00",x"00",x"00",x"00",x"0C",x"10",x"A8", -- 0x1478
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40", -- 0x1480
		x"BC",x"7F",x"F7",x"D7",x"B5",x"F7",x"FF",x"F7", -- 0x1488
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"42", -- 0x1490
		x"B9",x"FE",x"FA",x"7A",x"46",x"7E",x"7F",x"FF", -- 0x1498
		x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14A8
		x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x14B8
		x"55",x"5A",x"6B",x"A9",x"CB",x"36",x"11",x"2C", -- 0x14C0
		x"8A",x"82",x"C4",x"E3",x"F3",x"F8",x"F8",x"FC", -- 0x14C8
		x"55",x"8E",x"E5",x"22",x"D6",x"2D",x"03",x"D4", -- 0x14D0
		x"AA",x"91",x"EA",x"86",x"31",x"B2",x"AB",x"DA", -- 0x14D8
		x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"CF", -- 0x14E0
		x"CF",x"FF",x"83",x"FF",x"E7",x"E7",x"E7",x"E7", -- 0x14E8
		x"51",x"0A",x"29",x"90",x"84",x"CB",x"C5",x"E4", -- 0x14F0
		x"F0",x"F3",x"F0",x"F8",x"F9",x"FC",x"FC",x"FC", -- 0x14F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00", -- 0x1500
		x"7D",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1508
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00", -- 0x1510
		x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1520
		x"FF",x"00",x"FB",x"00",x"00",x"00",x"00",x"00", -- 0x1528
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1530
		x"FF",x"00",x"EF",x"00",x"00",x"00",x"00",x"00", -- 0x1538
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1540
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1548
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1550
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1558
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00", -- 0x1560
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1568
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00", -- 0x1570
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1578
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1580
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1588
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1590
		x"00",x"00",x"3E",x"7E",x"6E",x"C6",x"EE",x"FE", -- 0x1598
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15A8
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E8
		x"DE",x"DE",x"DE",x"DE",x"DE",x"DE",x"DE",x"DE", -- 0x15F0
		x"DE",x"DF",x"DF",x"DF",x"DF",x"FF",x"FF",x"FF", -- 0x15F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"BE",x"00", -- 0x1600
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1608
		x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"C0",x"7B", -- 0x1610
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1618
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1620
		x"3F",x"C0",x"2F",x"00",x"00",x"00",x"00",x"00", -- 0x1628
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1630
		x"FF",x"00",x"BE",x"00",x"00",x"00",x"00",x"00", -- 0x1638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1640
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1658
		x"8F",x"60",x"F6",x"33",x"11",x"00",x"00",x"00", -- 0x1660
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1668
		x"FF",x"07",x"73",x"1B",x"0B",x"18",x"00",x"00", -- 0x1670
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1678
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1680
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1688
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1690
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1698
		x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00", -- 0x16A0
		x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"00", -- 0x16A8
		x"FF",x"FF",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x16B0
		x"00",x"00",x"00",x"00",x"00",x"0C",x"10",x"A8", -- 0x16B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16D8
		x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x16E0
		x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x16E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x16F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"BB",x"40", -- 0x1700
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80", -- 0x1708
		x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"EF",x"00", -- 0x1710
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1718
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1720
		x"00",x"EF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1728
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1730
		x"00",x"BE",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1738
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1740
		x"FF",x"FF",x"FF",x"00",x"EF",x"01",x"00",x"00", -- 0x1748
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1750
		x"FF",x"FF",x"FF",x"FF",x"03",x"BD",x"01",x"00", -- 0x1758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1760
		x"00",x"00",x"00",x"00",x"00",x"10",x"20",x"21", -- 0x1768
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1770
		x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00", -- 0x1778
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1798
		x"FF",x"FF",x"FF",x"FF",x"FC",x"00",x"00",x"00", -- 0x17A0
		x"00",x"00",x"00",x"00",x"00",x"10",x"20",x"21", -- 0x17A8
		x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00", -- 0x17B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00", -- 0x17B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17C0
		x"FF",x"FE",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0", -- 0x17C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"E0", -- 0x17D0
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17D8
		x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",x"FE",x"FF", -- 0x17E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x17F0
		x"E0",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1800
		x"00",x"00",x"00",x"FF",x"00",x"FF",x"FF",x"FF", -- 0x1808
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1810
		x"00",x"00",x"00",x"80",x"7F",x"80",x"FF",x"DE", -- 0x1818
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1820
		x"00",x"FF",x"01",x"FC",x"FF",x"FF",x"FF",x"FF", -- 0x1828
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1830
		x"00",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF", -- 0x1838
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1840
		x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1848
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1850
		x"FF",x"80",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1858
		x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"C0", -- 0x1860
		x"FF",x"FF",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1868
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1870
		x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1878
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1880
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC", -- 0x1888
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1890
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1898
		x"80",x"C0",x"B8",x"C0",x"C0",x"E0",x"C0",x"90", -- 0x18A0
		x"30",x"70",x"C0",x"F7",x"31",x"36",x"60",x"8F", -- 0x18A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B0
		x"00",x"00",x"38",x"1B",x"0B",x"73",x"07",x"FF", -- 0x18B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
		x"FE",x"FE",x"CE",x"86",x"86",x"CE",x"7E",x"B8", -- 0x18E0
		x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E8
		x"FE",x"FE",x"E6",x"A6",x"A6",x"9E",x"9E",x"F9", -- 0x18F0
		x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1900
		x"FF",x"FF",x"FF",x"03",x"00",x"00",x"00",x"00", -- 0x1908
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1910
		x"FF",x"FF",x"FF",x"FF",x"0F",x"00",x"00",x"00", -- 0x1918
		x"00",x"00",x"00",x"F8",x"FC",x"0E",x"07",x"03", -- 0x1920
		x"C1",x"E0",x"70",x"38",x"18",x"18",x"18",x"18", -- 0x1928
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x1930
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x1938
		x"18",x"18",x"18",x"18",x"38",x"70",x"E0",x"C1", -- 0x1940
		x"03",x"07",x"0E",x"FC",x"F8",x"00",x"00",x"00", -- 0x1948
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x1950
		x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1958
		x"00",x"00",x"07",x"FC",x"03",x"FF",x"FF",x"FF", -- 0x1960
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1968
		x"00",x"1F",x"F0",x"0F",x"FF",x"FF",x"FF",x"FF", -- 0x1970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1978
		x"00",x"00",x"00",x"00",x"43",x"C3",x"00",x"00", -- 0x1980
		x"00",x"01",x"01",x"06",x"0B",x"08",x"0B",x"0B", -- 0x1988
		x"00",x"00",x"00",x"00",x"20",x"E1",x"00",x"00", -- 0x1990
		x"00",x"00",x"00",x"00",x"FE",x"0E",x"E0",x"2F", -- 0x1998
		x"08",x"0A",x"0B",x"89",x"8C",x"46",x"83",x"01", -- 0x19A0
		x"00",x"00",x"08",x"08",x"9F",x"FF",x"00",x"00", -- 0x19A8
		x"00",x"01",x"81",x"E0",x"FA",x"04",x"FA",x"02", -- 0x19B0
		x"0D",x"18",x"30",x"E7",x"CE",x"9C",x"38",x"70", -- 0x19B8
		x"03",x"FE",x"00",x"10",x"FF",x"00",x"00",x"00", -- 0x19C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19C8
		x"E4",x"04",x"48",x"F8",x"00",x"00",x"00",x"00", -- 0x19D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19D8
		x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00", -- 0x19E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19E8
		x"FE",x"AA",x"AA",x"6A",x"6E",x"BE",x"60",x"00", -- 0x19F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A00
		x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A10
		x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A18
		x"00",x"00",x"00",x"F0",x"F8",x"1C",x"0F",x"07", -- 0x1A20
		x"C3",x"E0",x"70",x"38",x"18",x"18",x"18",x"18", -- 0x1A28
		x"00",x"00",x"00",x"3F",x"7F",x"E0",x"C0",x"80", -- 0x1A30
		x"0F",x"1F",x"38",x"70",x"60",x"60",x"60",x"60", -- 0x1A38
		x"18",x"18",x"18",x"18",x"38",x"70",x"E0",x"C3", -- 0x1A40
		x"07",x"0F",x"1C",x"F8",x"F0",x"00",x"00",x"00", -- 0x1A48
		x"60",x"60",x"60",x"60",x"70",x"38",x"1F",x"0F", -- 0x1A50
		x"80",x"C0",x"E0",x"7F",x"3F",x"00",x"00",x"00", -- 0x1A58
		x"00",x"00",x"00",x"00",x"00",x"7F",x"80",x"7F", -- 0x1A60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A68
		x"00",x"00",x"00",x"00",x"7F",x"80",x"FF",x"FF", -- 0x1A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A78
		x"00",x"C7",x"00",x"00",x"00",x"FF",x"00",x"00", -- 0x1A80
		x"40",x"00",x"B8",x"82",x"84",x"80",x"A8",x"A8", -- 0x1A88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1A90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80", -- 0x1A98
		x"AA",x"AA",x"AE",x"A6",x"A6",x"B3",x"B8",x"BC", -- 0x1AA0
		x"3F",x"1E",x"00",x"00",x"0F",x"07",x"80",x"80", -- 0x1AA8
		x"80",x"C0",x"A0",x"70",x"00",x"F8",x"F8",x"03", -- 0x1AB0
		x"FE",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00", -- 0x1AB8
		x"20",x"00",x"9F",x"00",x"01",x"7F",x"80",x"00", -- 0x1AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AC8
		x"00",x"00",x"00",x"04",x"7F",x"80",x"00",x"00", -- 0x1AD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AD8
		x"02",x"04",x"04",x"01",x"00",x"01",x"01",x"02", -- 0x1AE0
		x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AE8
		x"00",x"18",x"20",x"50",x"A0",x"90",x"00",x"00", -- 0x1AF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1AF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"00", -- 0x1B00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x1B10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B18
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07", -- 0x1B20
		x"0E",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C", -- 0x1B28
		x"00",x"00",x"00",x"7F",x"FF",x"C0",x"80",x"00", -- 0x1B30
		x"0F",x"1F",x"38",x"70",x"60",x"60",x"60",x"60", -- 0x1B38
		x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0E", -- 0x1B40
		x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00", -- 0x1B48
		x"60",x"60",x"60",x"60",x"70",x"38",x"1F",x"0F", -- 0x1B50
		x"00",x"80",x"C0",x"FF",x"7F",x"00",x"00",x"00", -- 0x1B58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F", -- 0x1B60
		x"F0",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B68
		x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"80", -- 0x1B70
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B78
		x"00",x"FF",x"00",x"00",x"80",x"E0",x"38",x"02", -- 0x1B80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1B88
		x"00",x"FF",x"00",x"FF",x"08",x"28",x"28",x"28", -- 0x1B90
		x"2F",x"20",x"3F",x"23",x"21",x"90",x"14",x"14", -- 0x1B98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BA0
		x"00",x"00",x"E8",x"1A",x"E5",x"06",x"63",x"F3", -- 0x1BA8
		x"14",x"14",x"16",x"50",x"28",x"78",x"F8",x"F8", -- 0x1BB0
		x"3B",x"3B",x"3B",x"25",x"30",x"65",x"F3",x"07", -- 0x1BB8
		x"78",x"3C",x"1F",x"0F",x"00",x"04",x"FF",x"00", -- 0x1BC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BC8
		x"00",x"03",x"FF",x"FF",x"00",x"10",x"FF",x"00", -- 0x1BD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1BD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1ED8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x1FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
