-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_N2 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_N2 is


	type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0000
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0008
		x"BF",x"FF",x"BD",x"E3",x"F0",x"F1",x"9B",x"2F", -- 0x0010
		x"BD",x"EF",x"BD",x"EF",x"BD",x"EF",x"BD",x"EF", -- 0x0018
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x0020
		x"AD",x"FF",x"F8",x"FF",x"78",x"FF",x"78",x"DD", -- 0x0028
		x"78",x"DD",x"78",x"1D",x"F0",x"D1",x"0F",x"1D", -- 0x0030
		x"78",x"DD",x"78",x"DD",x"78",x"97",x"E3",x"E9", -- 0x0038
		x"BD",x"EF",x"BD",x"EF",x"BD",x"EF",x"BD",x"E3", -- 0x0040
		x"F0",x"F1",x"9B",x"2F",x"BF",x"FF",x"FF",x"FF", -- 0x0048
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0050
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
		x"0F",x"1F",x"78",x"DD",x"78",x"DD",x"78",x"1D", -- 0x0060
		x"F0",x"D1",x"0F",x"1D",x"78",x"DD",x"78",x"DD", -- 0x0068
		x"78",x"FF",x"F8",x"FF",x"AD",x"FF",x"DF",x"FF", -- 0x0070
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0078
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0080
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0088
		x"FF",x"FF",x"BF",x"EF",x"97",x"E3",x"78",x"79", -- 0x0090
		x"59",x"2F",x"9B",x"EF",x"9F",x"EF",x"9F",x"EF", -- 0x0098
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00A0
		x"DF",x"FF",x"8F",x"FF",x"AD",x"FF",x"2D",x"FF", -- 0x00A8
		x"2D",x"DD",x"2D",x"DD",x"F0",x"1D",x"F0",x"D1", -- 0x00B0
		x"3C",x"1D",x"3C",x"DD",x"78",x"95",x"F0",x"E1", -- 0x00B8
		x"9F",x"EF",x"9F",x"EF",x"9F",x"EF",x"97",x"E3", -- 0x00C0
		x"78",x"79",x"59",x"2F",x"BB",x"FF",x"FF",x"FF", -- 0x00C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00D8
		x"3F",x"9F",x"3C",x"DD",x"3C",x"DD",x"78",x"1D", -- 0x00E0
		x"F0",x"D1",x"0F",x"1D",x"3C",x"DD",x"3C",x"DD", -- 0x00E8
		x"3C",x"FF",x"BC",x"FF",x"AD",x"FF",x"DF",x"FF", -- 0x00F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x00F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0100
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0108
		x"FF",x"FF",x"BF",x"EF",x"5B",x"E3",x"1E",x"79", -- 0x0110
		x"1F",x"2F",x"BD",x"EF",x"BD",x"EF",x"BD",x"EF", -- 0x0118
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0120
		x"DF",x"FF",x"AD",x"FF",x"BC",x"FF",x"3C",x"FF", -- 0x0128
		x"3C",x"DD",x"3C",x"DD",x"F0",x"1D",x"F0",x"D1", -- 0x0130
		x"3C",x"1D",x"3C",x"DD",x"7B",x"9D",x"F0",x"E1", -- 0x0138
		x"BD",x"EF",x"BD",x"EF",x"BD",x"EF",x"79",x"E3", -- 0x0140
		x"1E",x"79",x"1B",x"2F",x"BF",x"FF",x"FF",x"FF", -- 0x0148
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0150
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0158
		x"0F",x"1F",x"3C",x"DD",x"3C",x"DD",x"78",x"1D", -- 0x0160
		x"F0",x"D1",x"0F",x"1D",x"3C",x"DD",x"3C",x"DD", -- 0x0168
		x"3C",x"FF",x"BC",x"FF",x"AD",x"FF",x"DF",x"FF", -- 0x0170
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0178
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0180
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0188
		x"BF",x"EF",x"1F",x"E3",x"2D",x"0F",x"5B",x"3F", -- 0x0190
		x"9F",x"EF",x"9F",x"EF",x"9F",x"EF",x"9F",x"EF", -- 0x0198
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x01A0
		x"8F",x"FF",x"8F",x"FF",x"1E",x"FF",x"1E",x"DD", -- 0x01A8
		x"1E",x"DD",x"1E",x"D1",x"0F",x"1D",x"0F",x"1D", -- 0x01B0
		x"0F",x"DD",x"1E",x"DD",x"3C",x"F1",x"0F",x"3C", -- 0x01B8
		x"9F",x"EF",x"9F",x"EF",x"1F",x"E3",x"2D",x"0F", -- 0x01C0
		x"5B",x"3F",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01D8
		x"3F",x"9F",x"0F",x"DD",x"1E",x"D1",x"0F",x"1D", -- 0x01E0
		x"0F",x"1D",x"0F",x"DD",x"1E",x"DD",x"0F",x"FF", -- 0x01E8
		x"8F",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x01F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0200
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0208
		x"FF",x"FF",x"BF",x"FF",x"9F",x"F3",x"1E",x"F0", -- 0x0210
		x"BD",x"2F",x"BD",x"EF",x"BD",x"EF",x"BD",x"EF", -- 0x0218
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0220
		x"FF",x"FF",x"DF",x"FF",x"AD",x"FF",x"BC",x"FF", -- 0x0228
		x"3C",x"DD",x"3C",x"DD",x"F0",x"95",x"F0",x"1D", -- 0x0230
		x"78",x"1D",x"78",x"DD",x"7B",x"DB",x"78",x"E1", -- 0x0238
		x"BD",x"EF",x"BD",x"EF",x"BD",x"EF",x"9F",x"F3", -- 0x0240
		x"1E",x"F0",x"BD",x"2E",x"FB",x"FF",x"FF",x"FF", -- 0x0248
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0250
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0258
		x"0F",x"1F",x"3C",x"DD",x"3C",x"DD",x"F0",x"95", -- 0x0260
		x"F0",x"1D",x"3C",x"1D",x"3C",x"DD",x"3C",x"DD", -- 0x0268
		x"3C",x"FF",x"AD",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x0270
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0278
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0280
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0288
		x"FF",x"FF",x"3F",x"EF",x"97",x"E3",x"09",x"0F", -- 0x0290
		x"1B",x"3F",x"9F",x"EF",x"9F",x"EF",x"9F",x"EF", -- 0x0298
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02A0
		x"FF",x"FF",x"DF",x"FF",x"8F",x"FF",x"0F",x"FF", -- 0x02A8
		x"0F",x"DD",x"0F",x"D5",x"0F",x"59",x"0F",x"1D", -- 0x02B0
		x"0F",x"DD",x"0F",x"DD",x"0F",x"D1",x"0F",x"2D", -- 0x02B8
		x"1F",x"EF",x"97",x"E3",x"09",x"0F",x"1B",x"3F", -- 0x02C0
		x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02D8
		x"3F",x"9F",x"0F",x"59",x"0F",x"1D",x"0F",x"DD", -- 0x02E0
		x"0F",x"DD",x"0F",x"DD",x"8F",x"FF",x"DF",x"FF", -- 0x02E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0300
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0308
		x"FF",x"FF",x"FF",x"FF",x"FB",x"FF",x"F9",x"F3", -- 0x0310
		x"1E",x"F0",x"BD",x"2F",x"BD",x"EF",x"BD",x"EF", -- 0x0318
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0320
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x0328
		x"AD",x"FF",x"3C",x"DD",x"3C",x"DD",x"3C",x"DD", -- 0x0330
		x"F0",x"D1",x"78",x"95",x"7B",x"DB",x"78",x"E1", -- 0x0338
		x"BD",x"EF",x"BD",x"EF",x"BD",x"F3",x"1E",x"F0", -- 0x0340
		x"BD",x"2E",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0348
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0350
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0358
		x"0F",x"1D",x"3C",x"DD",x"3C",x"DD",x"F0",x"95", -- 0x0360
		x"F0",x"1D",x"3C",x"5D",x"34",x"DD",x"BC",x"FF", -- 0x0368
		x"AD",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0370
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0378
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0380
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0388
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x0390
		x"F0",x"FF",x"F0",x"F7",x"FF",x"F0",x"FF",x"F8", -- 0x0398
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F3",x"FF", -- 0x03B0
		x"FB",x"FF",x"FB",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x03B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"F4", -- 0x03D0
		x"F7",x"F8",x"F7",x"FB",x"F0",x"F3",x"F0",x"F4", -- 0x03D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x03E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F3",x"FF", -- 0x03F0
		x"F3",x"FF",x"FB",x"FF",x"FB",x"FF",x"F3",x"FF", -- 0x03F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0400
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x0408
		x"DF",x"EF",x"CF",x"EF",x"CF",x"CB",x"E9",x"0F", -- 0x0410
		x"CC",x"EF",x"CD",x"EF",x"CF",x"EF",x"CF",x"EF", -- 0x0418
		x"FF",x"FF",x"FF",x"FF",x"FB",x"FF",x"1F",x"FF", -- 0x0420
		x"3D",x"FF",x"3D",x"FF",x"3D",x"FF",x"3D",x"FF", -- 0x0428
		x"3C",x"3F",x"0F",x"BF",x"0F",x"7F",x"1F",x"FF", -- 0x0430
		x"3D",x"FF",x"3D",x"FF",x"3C",x"B7",x"6F",x"5B", -- 0x0438
		x"CF",x"EF",x"CF",x"EF",x"CF",x"EB",x"E9",x"0F", -- 0x0440
		x"CC",x"8F",x"CD",x"EF",x"DF",x"EF",x"FF",x"EF", -- 0x0448
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0450
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0458
		x"0F",x"3F",x"1F",x"FF",x"3D",x"FF",x"3D",x"FF", -- 0x0460
		x"3C",x"7F",x"0F",x"BF",x"0F",x"3B",x"1F",x"FF", -- 0x0468
		x"3D",x"FF",x"3D",x"FF",x"3D",x"FF",x"3D",x"FF", -- 0x0470
		x"1F",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0480
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0488
		x"FF",x"EF",x"FF",x"AF",x"FF",x"8F",x"FF",x"1B", -- 0x0490
		x"FE",x"3F",x"FF",x"BF",x"FF",x"BF",x"FF",x"BF", -- 0x0498
		x"FF",x"FF",x"BF",x"FF",x"BF",x"FF",x"3F",x"FF", -- 0x04A0
		x"3F",x"FF",x"3F",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x04A8
		x"1F",x"FF",x"0F",x"FF",x"02",x"FF",x"3F",x"FF", -- 0x04B0
		x"3F",x"FF",x"3F",x"FF",x"0F",x"FF",x"4F",x"7F", -- 0x04B8
		x"FF",x"BF",x"FF",x"BF",x"FE",x"3F",x"FF",x"1F", -- 0x04C0
		x"FF",x"8B",x"FF",x"AF",x"FF",x"FF",x"FF",x"FF", -- 0x04C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04D8
		x"07",x"FF",x"3B",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x04E0
		x"0F",x"FF",x"0F",x"FF",x"17",x"FF",x"3B",x"FF", -- 0x04E8
		x"3F",x"FF",x"3F",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x04F0
		x"BF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x04F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"9F",x"FF",x"9F", -- 0x0500
		x"FF",x"9F",x"FF",x"BD",x"FF",x"AD",x"FF",x"AD", -- 0x0508
		x"DF",x"96",x"CF",x"E1",x"EF",x"3C",x"FF",x"0F", -- 0x0510
		x"FF",x"8F",x"FF",x"AD",x"8F",x"3C",x"BC",x"C3", -- 0x0518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0520
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0528
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"A7",x"FF", -- 0x0530
		x"5A",x"FF",x"8F",x"7B",x"CF",x"7F",x"FE",x"FF", -- 0x0538
		x"8F",x"1E",x"FF",x"AD",x"FF",x"BC",x"FF",x"1E", -- 0x0540
		x"EF",x"69",x"DF",x"C3",x"CF",x"1E",x"FF",x"AD", -- 0x0548
		x"FF",x"AD",x"FF",x"BD",x"FF",x"9F",x"FF",x"9F", -- 0x0550
		x"FF",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0558
		x"FE",x"FF",x"FC",x"F7",x"BC",x"7B",x"87",x"FF", -- 0x0560
		x"2F",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0568
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0570
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0578
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"EF", -- 0x0580
		x"FF",x"EF",x"FF",x"EF",x"FF",x"EF",x"FF",x"EF", -- 0x0588
		x"FF",x"EF",x"FF",x"DE",x"FF",x"CE",x"FF",x"CF", -- 0x0590
		x"FF",x"CD",x"FF",x"EF",x"FF",x"AD",x"FF",x"8F", -- 0x0598
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"FF", -- 0x05A8
		x"FB",x"FF",x"F0",x"FF",x"3B",x"FF",x"3F",x"FF", -- 0x05B0
		x"7B",x"FF",x"FB",x"FF",x"F3",x"FF",x"7B",x"FF", -- 0x05B8
		x"FF",x"8F",x"FF",x"EF",x"FF",x"CD",x"FF",x"CF", -- 0x05C0
		x"FF",x"CF",x"FF",x"FE",x"FF",x"EE",x"FF",x"EF", -- 0x05C8
		x"FF",x"EF",x"FF",x"EF",x"FF",x"EF",x"FF",x"EF", -- 0x05D0
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05D8
		x"7B",x"FF",x"FB",x"FF",x"7B",x"FF",x"7B",x"FF", -- 0x05E0
		x"F3",x"FF",x"F0",x"FF",x"BB",x"FF",x"BF",x"FF", -- 0x05E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0600
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0608
		x"FF",x"EF",x"FF",x"4F",x"FF",x"0F",x"EF",x"0F", -- 0x0610
		x"ED",x"37",x"FF",x"7F",x"FF",x"7F",x"FF",x"7F", -- 0x0618
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"9F",x"FF", -- 0x0620
		x"9F",x"FF",x"9F",x"FF",x"1F",x"FF",x"1F",x"FF", -- 0x0628
		x"1E",x"7F",x"0F",x"BF",x"0F",x"77",x"1F",x"FF", -- 0x0630
		x"1F",x"FF",x"1F",x"FF",x"1E",x"7F",x"6F",x"3F", -- 0x0638
		x"FF",x"7F",x"FF",x"7F",x"ED",x"3F",x"EF",x"0F", -- 0x0640
		x"FF",x"07",x"FF",x"4F",x"FF",x"FF",x"FF",x"FF", -- 0x0648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0658
		x"0F",x"77",x"1F",x"FF",x"1F",x"FF",x"1F",x"FF", -- 0x0660
		x"1E",x"7F",x"0F",x"BF",x"0F",x"77",x"1F",x"FF", -- 0x0668
		x"1F",x"FF",x"9F",x"FF",x"9F",x"FF",x"9F",x"FF", -- 0x0670
		x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x0680
		x"FF",x"FE",x"FF",x"FE",x"FF",x"FE",x"FF",x"FE", -- 0x0688
		x"FF",x"CE",x"FF",x"9E",x"FF",x"CE",x"FF",x"AF", -- 0x0690
		x"FF",x"9E",x"EF",x"3E",x"FF",x"DE",x"FF",x"8F", -- 0x0698
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06A8
		x"7F",x"FF",x"B7",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x06B0
		x"FF",x"FF",x"FF",x"FF",x"3F",x"FF",x"B7",x"FF", -- 0x06B8
		x"FF",x"DE",x"EF",x"2E",x"FF",x"8F",x"FF",x"BE", -- 0x06C0
		x"FF",x"DE",x"FF",x"9E",x"FF",x"CE",x"FF",x"EE", -- 0x06C8
		x"FF",x"EF",x"FF",x"FE",x"FF",x"FE",x"FF",x"EF", -- 0x06D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06D8
		x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06E0
		x"7F",x"FF",x"B7",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x06E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"DF", -- 0x0700
		x"FF",x"CF",x"FF",x"CF",x"FF",x"CF",x"FF",x"CF", -- 0x0708
		x"FF",x"CF",x"FF",x"CF",x"FF",x"8F",x"FF",x"0F", -- 0x0710
		x"FF",x"06",x"FF",x"CD",x"FF",x"0F",x"EF",x"0F", -- 0x0718
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0720
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F", -- 0x0728
		x"7F",x"7F",x"0F",x"F1",x"0F",x"77",x"3F",x"7F", -- 0x0730
		x"77",x"7F",x"3F",x"7F",x"3F",x"7F",x"3F",x"7F", -- 0x0738
		x"FF",x"07",x"FF",x"CC",x"FF",x"0F",x"FF",x"0F", -- 0x0740
		x"FF",x"8B",x"FF",x"CE",x"FF",x"CF",x"FF",x"CF", -- 0x0748
		x"FF",x"CF",x"FF",x"CF",x"FF",x"CF",x"FF",x"CF", -- 0x0750
		x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0758
		x"37",x"7F",x"3F",x"7F",x"7F",x"7F",x"3F",x"7F", -- 0x0760
		x"0F",x"7F",x"0F",x"F1",x"7F",x"77",x"7F",x"7F", -- 0x0768
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"FB", -- 0x0788
		x"FF",x"7B",x"FF",x"38",x"FF",x"EB",x"FF",x"FB", -- 0x0790
		x"FF",x"FB",x"FF",x"FB",x"FF",x"FB",x"FF",x"FB", -- 0x0798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"FF", -- 0x07A0
		x"7B",x"FF",x"7B",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x07A8
		x"F3",x"FF",x"97",x"FF",x"F1",x"FF",x"1F",x"FF", -- 0x07B0
		x"B7",x"FF",x"F3",x"FF",x"D3",x"FF",x"A7",x"FF", -- 0x07B8
		x"FF",x"FB",x"FF",x"FB",x"FF",x"FB",x"FF",x"FB", -- 0x07C0
		x"FF",x"EB",x"FF",x"78",x"FF",x"F3",x"FF",x"BB", -- 0x07C8
		x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07D8
		x"1F",x"FF",x"B7",x"FF",x"F3",x"FF",x"D3",x"FF", -- 0x07E0
		x"F1",x"FF",x"97",x"FF",x"3F",x"FF",x"F3",x"FF", -- 0x07E8
		x"F3",x"FF",x"7B",x"FF",x"7B",x"FF",x"BF",x"FF", -- 0x07F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x07F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0800
		x"FF",x"FF",x"FF",x"FF",x"FE",x"7F",x"DE",x"F7", -- 0x0808
		x"CF",x"E7",x"CE",x"69",x"CD",x"16",x"FE",x"4F", -- 0x0810
		x"FE",x"F7",x"FE",x"F7",x"FE",x"F7",x"FE",x"F7", -- 0x0818
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x0820
		x"BD",x"FF",x"F9",x"FF",x"79",x"FF",x"79",x"FF", -- 0x0828
		x"F1",x"FF",x"E1",x"FF",x"F0",x"7F",x"0F",x"7F", -- 0x0830
		x"F1",x"FF",x"F1",x"FF",x"69",x"FF",x"F6",x"7F", -- 0x0838
		x"FE",x"F7",x"FE",x"F7",x"FE",x"F7",x"FE",x"C7", -- 0x0840
		x"FC",x"B4",x"FC",x"E1",x"FC",x"6F",x"EF",x"FF", -- 0x0848
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0850
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0858
		x"0F",x"FF",x"97",x"FF",x"F1",x"FF",x"E1",x"7F", -- 0x0860
		x"F0",x"7F",x"0F",x"FF",x"1F",x"FF",x"79",x"FF", -- 0x0868
		x"F9",x"FF",x"F9",x"FF",x"BD",x"FF",x"DF",x"FF", -- 0x0870
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0878
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0880
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0888
		x"7F",x"FD",x"B5",x"F9",x"78",x"97",x"0F",x"78", -- 0x0890
		x"7F",x"09",x"F7",x"B9",x"F7",x"F9",x"F7",x"F9", -- 0x0898
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08B8
		x"F7",x"F9",x"F7",x"F9",x"F7",x"F9",x"F7",x"96", -- 0x08C0
		x"78",x"78",x"E1",x"19",x"1F",x"B9",x"7F",x"DF", -- 0x08C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x08F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0900
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0908
		x"5E",x"6F",x"F0",x"2F",x"0F",x"C3",x"4D",x"4E", -- 0x0910
		x"7F",x"EE",x"7F",x"EE",x"7F",x"EF",x"7F",x"EF", -- 0x0918
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0920
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x0928
		x"B7",x"FF",x"F3",x"FF",x"5B",x"FF",x"3C",x"FF", -- 0x0930
		x"37",x"FF",x"F3",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x0938
		x"7F",x"EF",x"7F",x"EF",x"7F",x"EF",x"7F",x"EF", -- 0x0940
		x"5E",x"E5",x"3C",x"0F",x"87",x"2E",x"4D",x"6E", -- 0x0948
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0950
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0958
		x"F3",x"FF",x"F3",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x0960
		x"B4",x"FF",x"D3",x"FF",x"37",x"FF",x"B7",x"FF", -- 0x0968
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0978
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0980
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0988
		x"DB",x"FF",x"F9",x"6B",x"78",x"D3",x"B9",x"2F", -- 0x0990
		x"BD",x"EF",x"BD",x"EF",x"BD",x"EF",x"BD",x"EF", -- 0x0998
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x09A0
		x"8F",x"FF",x"AD",x"FF",x"2D",x"FF",x"2D",x"FF", -- 0x09A8
		x"2D",x"BB",x"78",x"3B",x"0F",x"3B",x"0F",x"3B", -- 0x09B0
		x"0F",x"BB",x"2D",x"FF",x"78",x"3F",x"3F",x"97", -- 0x09B8
		x"BD",x"EF",x"BD",x"EF",x"BD",x"6B",x"78",x"D3", -- 0x09C0
		x"B9",x"2F",x"DB",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x09C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09D8
		x"0F",x"3F",x"2D",x"BB",x"F0",x"3B",x"0F",x"3B", -- 0x09E0
		x"0F",x"3B",x"0F",x"BB",x"2D",x"FF",x"2D",x"FF", -- 0x09E8
		x"AD",x"FF",x"8F",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x09F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A00
		x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"FC",x"FF", -- 0x0A08
		x"BC",x"F9",x"9E",x"F0",x"CC",x"8F",x"FC",x"FF", -- 0x0A10
		x"FC",x"FF",x"FC",x"FF",x"FC",x"FF",x"FC",x"FF", -- 0x0A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x0A20
		x"9F",x"FF",x"DB",x"FF",x"5B",x"FF",x"5B",x"FF", -- 0x0A28
		x"D3",x"FF",x"F8",x"7F",x"F0",x"7F",x"0F",x"7F", -- 0x0A30
		x"D3",x"FF",x"D3",x"FF",x"B4",x"7F",x"7E",x"B7", -- 0x0A38
		x"FC",x"FF",x"FC",x"FF",x"FC",x"FF",x"FC",x"FF", -- 0x0A40
		x"FC",x"BC",x"F8",x"F0",x"C9",x"9F",x"FD",x"FF", -- 0x0A48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A58
		x"0F",x"7F",x"97",x"FF",x"D3",x"FF",x"F0",x"F7", -- 0x0A60
		x"F0",x"F7",x"8F",x"7F",x"5B",x"FF",x"5B",x"FF", -- 0x0A68
		x"DB",x"FF",x"DB",x"FF",x"9F",x"FF",x"DF",x"FF", -- 0x0A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0A90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x0A98
		x"FF",x"FF",x"FF",x"BF",x"FF",x"9F",x"FF",x"DB", -- 0x0AA0
		x"FF",x"F9",x"FF",x"E9",x"FF",x"E9",x"CE",x"78", -- 0x0AA8
		x"CF",x"F0",x"CF",x"78",x"EF",x"0F",x"FF",x"8F", -- 0x0AB0
		x"FF",x"F8",x"FF",x"F8",x"0F",x"78",x"78",x"87", -- 0x0AB8
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0AD8
		x"3C",x"C3",x"0F",x"1E",x"FF",x"F8",x"FF",x"F8", -- 0x0AE0
		x"FF",x"E9",x"EF",x"1E",x"CF",x"78",x"CE",x"C3", -- 0x0AE8
		x"CF",x"1E",x"FF",x"F8",x"FF",x"E9",x"FF",x"E9", -- 0x0AF0
		x"FF",x"DB",x"FF",x"9F",x"FF",x"BF",x"FF",x"FF", -- 0x0AF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"CF", -- 0x0B18
		x"FF",x"BF",x"FF",x"5B",x"FF",x"79",x"FF",x"79", -- 0x0B20
		x"FF",x"69",x"FF",x"78",x"FF",x"78",x"CF",x"78", -- 0x0B28
		x"9A",x"F0",x"8F",x"1E",x"CF",x"0F",x"FF",x"78", -- 0x0B30
		x"FF",x"78",x"FF",x"78",x"0F",x"78",x"F0",x"D2", -- 0x0B38
		x"FF",x"CF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x0B40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B58
		x"78",x"87",x"0F",x"1E",x"FF",x"3C",x"FF",x"78", -- 0x0B60
		x"FF",x"78",x"CF",x"78",x"8F",x"F0",x"9A",x"87", -- 0x0B68
		x"CF",x"1E",x"FF",x"78",x"FF",x"78",x"FF",x"69", -- 0x0B70
		x"FF",x"79",x"FF",x"79",x"FF",x"5B",x"FF",x"BF", -- 0x0B78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0B88
		x"FF",x"FF",x"DF",x"FF",x"CF",x"AF",x"BC",x"F1", -- 0x0B90
		x"CD",x"AF",x"CF",x"EF",x"CF",x"EF",x"CF",x"EF", -- 0x0B98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BA0
		x"FF",x"FF",x"DF",x"FF",x"CF",x"FF",x"AD",x"FF", -- 0x0BA8
		x"AD",x"FF",x"2D",x"BB",x"2D",x"BB",x"F0",x"3B", -- 0x0BB0
		x"0F",x"3B",x"0F",x"BB",x"3C",x"3F",x"7B",x"97", -- 0x0BB8
		x"CF",x"EF",x"CF",x"EF",x"CF",x"AF",x"BC",x"F1", -- 0x0BC0
		x"CD",x"AF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BD8
		x"0F",x"3F",x"0F",x"BB",x"2D",x"BB",x"F0",x"3B", -- 0x0BE0
		x"0F",x"3B",x"0F",x"BB",x"AD",x"FF",x"AD",x"FF", -- 0x0BE8
		x"CF",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0BF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C10
		x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x0C18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C30
		x"FF",x"FF",x"FB",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x0C38
		x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"F7",x"FE", -- 0x0C40
		x"F0",x"F0",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x0C48
		x"F7",x"FE",x"F0",x"F0",x"FF",x"FF",x"F0",x"F0", -- 0x0C50
		x"F0",x"F0",x"F7",x"FE",x"F0",x"F0",x"FF",x"FF", -- 0x0C58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0C88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F1",x"F8", -- 0x0C90
		x"F7",x"F8",x"F7",x"FB",x"F0",x"F3",x"F0",x"F3", -- 0x0C98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F3",x"FF", -- 0x0CB0
		x"F3",x"FF",x"FB",x"FF",x"FB",x"FF",x"FB",x"FF", -- 0x0CB8
		x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"F7",x"FE", -- 0x0CC0
		x"F0",x"F0",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x0CC8
		x"F7",x"FE",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x0CD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0CF8
		x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"F7",x"FE", -- 0x0D00
		x"F0",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D38
		x"FC",x"F7",x"FB",x"FF",x"FB",x"FF",x"FB",x"FF", -- 0x0D40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FF", -- 0x0D50
		x"FB",x"FF",x"FB",x"FF",x"FC",x"F7",x"FF",x"FF", -- 0x0D58
		x"FF",x"F1",x"FF",x"FE",x"FF",x"FE",x"FF",x"FE", -- 0x0D60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x0D70
		x"FF",x"FE",x"FF",x"FE",x"FF",x"F1",x"FF",x"FF", -- 0x0D78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D80
		x"FF",x"7F",x"EF",x"97",x"FF",x"3F",x"FF",x"3F", -- 0x0D88
		x"FF",x"3F",x"FF",x"3F",x"EF",x"97",x"FF",x"7F", -- 0x0D90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D98
		x"9F",x"FF",x"9F",x"FF",x"9F",x"FF",x"1F",x"FF", -- 0x0DA0
		x"0F",x"FF",x"0F",x"FF",x"1F",x"FF",x"3C",x"7F", -- 0x0DA8
		x"6F",x"7F",x"1F",x"FF",x"0F",x"FF",x"0F",x"FF", -- 0x0DB0
		x"1F",x"FF",x"9F",x"FF",x"9F",x"FF",x"9F",x"FF", -- 0x0DB8
		x"FF",x"FF",x"FF",x"EE",x"FF",x"EE",x"FF",x"6F", -- 0x0DC0
		x"EF",x"97",x"CC",x"09",x"EE",x"4D",x"EE",x"4D", -- 0x0DC8
		x"EE",x"4D",x"EE",x"4D",x"EF",x"97",x"CC",x"09", -- 0x0DD0
		x"EE",x"66",x"FF",x"EE",x"FF",x"EE",x"FF",x"FF", -- 0x0DD8
		x"3F",x"FF",x"3F",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x0DE0
		x"D3",x"FF",x"3F",x"FF",x"5B",x"FF",x"E5",x"FF", -- 0x0DE8
		x"1F",x"FF",x"3F",x"FF",x"D3",x"FF",x"3F",x"FF", -- 0x0DF0
		x"3F",x"FF",x"3F",x"FF",x"3F",x"FF",x"77",x"FF", -- 0x0DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF", -- 0x0E08
		x"BD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DE", -- 0x0E48
		x"FF",x"DE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"B7",x"FF", -- 0x0E68
		x"B7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DE",x"FF",x"DE", -- 0x0E80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DE", -- 0x0E90
		x"FF",x"DE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E98
		x"FF",x"FF",x"FF",x"FF",x"B7",x"FF",x"B7",x"FF", -- 0x0EA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"B7",x"FF", -- 0x0EB0
		x"B7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BD",x"FF", -- 0x0EC8
		x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0ED8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DE", -- 0x0F08
		x"FF",x"DE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"B7",x"FF", -- 0x0F28
		x"B7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F30
		x"69",x"FF",x"69",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DE",x"FF",x"DE", -- 0x0F48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F58
		x"FF",x"FF",x"69",x"FF",x"69",x"FF",x"FF",x"FF", -- 0x0F60
		x"FF",x"FF",x"FF",x"FF",x"B7",x"FF",x"B7",x"FF", -- 0x0F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F78
		x"FF",x"FE",x"FF",x"DC",x"FF",x"30",x"EE",x"30", -- 0x0F80
		x"CC",x"70",x"DD",x"70",x"99",x"B8",x"99",x"DC", -- 0x0F88
		x"F0",x"F0",x"B8",x"E0",x"CC",x"C0",x"CC",x"22", -- 0x0F90
		x"EE",x"66",x"FF",x"00",x"FF",x"CC",x"FF",x"FF", -- 0x0F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA0
		x"FF",x"FF",x"FC",x"FF",x"F8",x"F3",x"F0",x"F0", -- 0x0FA8
		x"80",x"11",x"F3",x"DD",x"F1",x"FF",x"F1",x"BB", -- 0x0FB0
		x"F3",x"77",x"C0",x"FF",x"B3",x"FF",x"F7",x"FF", -- 0x0FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1000
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DE",x"F7", -- 0x1008
		x"F0",x"D3",x"0F",x"0F",x"0F",x"1D",x"CF",x"7F", -- 0x1010
		x"7F",x"FF",x"7F",x"FF",x"7F",x"FF",x"7F",x"FF", -- 0x1018
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1020
		x"FF",x"FF",x"DF",x"FF",x"8F",x"FF",x"8F",x"FF", -- 0x1028
		x"8F",x"FF",x"F0",x"F7",x"88",x"FF",x"89",x"FF", -- 0x1030
		x"8F",x"FF",x"8F",x"FF",x"8F",x"FF",x"8F",x"FF", -- 0x1038
		x"7F",x"FF",x"7F",x"FF",x"7F",x"FF",x"7F",x"FF", -- 0x1040
		x"DE",x"F7",x"F0",x"97",x"0F",x"0F",x"0F",x"1D", -- 0x1048
		x"CF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1050
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1058
		x"8F",x"FF",x"8F",x"FF",x"8F",x"FF",x"8F",x"FF", -- 0x1060
		x"8F",x"FF",x"8F",x"FF",x"F0",x"F7",x"88",x"FF", -- 0x1068
		x"89",x"FF",x"8F",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x1070
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1078
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1080
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x1088
		x"5E",x"ED",x"F0",x"E1",x"0F",x"6E",x"3F",x"EE", -- 0x1090
		x"7F",x"EE",x"7F",x"EF",x"3F",x"EF",x"3F",x"EF", -- 0x1098
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10A0
		x"FF",x"FF",x"FF",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x10A8
		x"D3",x"FF",x"3D",x"FF",x"33",x"FF",x"37",x"FF", -- 0x10B0
		x"3F",x"FF",x"3F",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x10B8
		x"3F",x"EF",x"3F",x"EF",x"7F",x"EF",x"7F",x"EF", -- 0x10C0
		x"3F",x"EF",x"0F",x"E7",x"F0",x"D2",x"4F",x"0E", -- 0x10C8
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10D8
		x"3F",x"FF",x"3F",x"FF",x"3F",x"FF",x"3F",x"FF", -- 0x10E0
		x"3F",x"FF",x"3F",x"FF",x"3D",x"FF",x"D3",x"FF", -- 0x10E8
		x"37",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x10F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1100
		x"7F",x"FF",x"7F",x"FF",x"7F",x"FF",x"3F",x"CF", -- 0x1108
		x"3E",x"CF",x"0F",x"1E",x"0F",x"4C",x"23",x"CD", -- 0x1110
		x"3F",x"CF",x"3F",x"CF",x"3F",x"CF",x"B7",x"CF", -- 0x1118
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1120
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1128
		x"FF",x"FF",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1130
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1138
		x"3F",x"CF",x"3F",x"CF",x"3F",x"CF",x"3F",x"CF", -- 0x1140
		x"3E",x"CF",x"0F",x"4F",x"0F",x"1E",x"23",x"CC", -- 0x1148
		x"3F",x"EF",x"7F",x"FF",x"7F",x"FF",x"7F",x"FF", -- 0x1150
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1158
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1160
		x"FF",x"FF",x"FF",x"FF",x"F3",x"FF",x"FF",x"FF", -- 0x1168
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1170
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1178
		x"FF",x"FF",x"CD",x"0F",x"CD",x"0F",x"CC",x"00", -- 0x1180
		x"CD",x"0E",x"CD",x"02",x"CD",x"0E",x"CC",x"00", -- 0x1188
		x"EE",x"1F",x"CD",x"19",x"CC",x"1F",x"CD",x"19", -- 0x1190
		x"CC",x"1F",x"EE",x"11",x"FF",x"FF",x"FF",x"FF", -- 0x1198
		x"FF",x"FF",x"0F",x"FF",x"0F",x"FF",x"09",x"FF", -- 0x11A0
		x"09",x"FF",x"0F",x"FF",x"0F",x"FF",x"00",x"FF", -- 0x11A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11B8
		x"FF",x"FF",x"FD",x"FF",x"FD",x"FF",x"FC",x"F0", -- 0x11C0
		x"FD",x"FE",x"FD",x"F2",x"FD",x"FE",x"FC",x"F0", -- 0x11C8
		x"FE",x"FF",x"FD",x"F9",x"FC",x"FF",x"FD",x"F9", -- 0x11D0
		x"FC",x"FF",x"FE",x"F1",x"FF",x"FF",x"FF",x"FF", -- 0x11D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF", -- 0x11E0
		x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"FF", -- 0x11E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1200
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"EE", -- 0x1208
		x"FF",x"EE",x"FF",x"EE",x"FF",x"EE",x"FF",x"EE", -- 0x1210
		x"FF",x"EE",x"FF",x"FF",x"FF",x"BC",x"FF",x"78", -- 0x1218
		x"FF",x"3F",x"EF",x"3F",x"EF",x"1F",x"EF",x"1F", -- 0x1220
		x"EF",x"1F",x"EF",x"0F",x"EF",x"0F",x"EF",x"0F", -- 0x1228
		x"78",x"F0",x"0F",x"0F",x"0F",x"0F",x"EE",x"00", -- 0x1230
		x"EF",x"0F",x"EF",x"0F",x"F0",x"C3",x"F0",x"F0", -- 0x1238
		x"FF",x"0F",x"FF",x"8F",x"FF",x"FF",x"FF",x"EE", -- 0x1240
		x"FF",x"EE",x"FF",x"EE",x"FF",x"EE",x"FF",x"EE", -- 0x1248
		x"FF",x"EE",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x1250
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1258
		x"0F",x"0F",x"0F",x"09",x"EE",x"07",x"EF",x"0F", -- 0x1260
		x"EF",x"0F",x"78",x"F0",x"0F",x"0F",x"0F",x"0F", -- 0x1268
		x"EE",x"00",x"EF",x"0F",x"EF",x"0F",x"EF",x"1F", -- 0x1270
		x"EF",x"1F",x"EF",x"1F",x"EF",x"3F",x"FF",x"3F", -- 0x1278
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1280
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1288
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1290
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"CF", -- 0x1298
		x"FF",x"FF",x"FF",x"BF",x"FF",x"1F",x"FF",x"1F", -- 0x12A0
		x"FF",x"1F",x"FF",x"0F",x"FF",x"0F",x"FF",x"0F", -- 0x12A8
		x"FF",x"0F",x"0F",x"1E",x"1E",x"E1",x"0F",x"0C", -- 0x12B0
		x"FF",x"03",x"FF",x"0F",x"0F",x"0F",x"0F",x"4B", -- 0x12B8
		x"FF",x"CD",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x12C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x12D8
		x"0F",x"0F",x"0F",x"0C",x"FF",x"03",x"FF",x"0F", -- 0x12E0
		x"0F",x"0F",x"78",x"E1",x"0F",x"1E",x"FF",x"03", -- 0x12E8
		x"FF",x"0F",x"FF",x"0F",x"FF",x"0F",x"FF",x"1F", -- 0x12F0
		x"FF",x"1F",x"FF",x"1F",x"FF",x"BF",x"FF",x"FF", -- 0x12F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1300
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1308
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1310
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1318
		x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"FF",x"CF", -- 0x1320
		x"FF",x"CF",x"FF",x"CF",x"FF",x"CF",x"FF",x"CF", -- 0x1328
		x"FF",x"CF",x"FF",x"0F",x"EF",x"0F",x"FF",x"04", -- 0x1330
		x"FF",x"CF",x"FF",x"CF",x"CF",x"2D",x"8F",x"0F", -- 0x1338
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1340
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1348
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1350
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1358
		x"8F",x"0F",x"CD",x"0E",x"FF",x"CD",x"FF",x"CF", -- 0x1360
		x"FF",x"0F",x"EF",x"0F",x"FF",x"07",x"FF",x"CC", -- 0x1368
		x"FF",x"CF",x"FF",x"CF",x"FF",x"CF",x"FF",x"CF", -- 0x1370
		x"FF",x"CF",x"FF",x"CF",x"FF",x"FF",x"FF",x"FF", -- 0x1378
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1380
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1388
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1390
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1398
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x13F8
		x"78",x"F0",x"3C",x"F0",x"0F",x"0F",x"0F",x"0F", -- 0x1400
		x"1E",x"1F",x"1E",x"2F",x"1E",x"4F",x"1E",x"5F", -- 0x1408
		x"1E",x"5F",x"1E",x"2F",x"1E",x"1F",x"1E",x"0F", -- 0x1410
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1418
		x"F0",x"F0",x"F0",x"F0",x"0F",x"3C",x"0F",x"3C", -- 0x1420
		x"CF",x"3C",x"2F",x"3C",x"9F",x"3C",x"5F",x"3C", -- 0x1428
		x"5F",x"3C",x"2F",x"3C",x"CF",x"3C",x"0F",x"3C", -- 0x1430
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x1438
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1440
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1448
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1450
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1458
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x1460
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x1468
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x1470
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x1478
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1480
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1488
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1490
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x1498
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x14A0
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x14A8
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x14B0
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x14B8
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x14C0
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x14C8
		x"1E",x"0F",x"1E",x"0F",x"1E",x"0F",x"1E",x"0F", -- 0x14D0
		x"1E",x"0F",x"1E",x"F0",x"0F",x"0F",x"0F",x"0F", -- 0x14D8
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x14E0
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x14E8
		x"0F",x"3C",x"0F",x"3C",x"0F",x"3C",x"0F",x"3C", -- 0x14F0
		x"0F",x"3C",x"F0",x"3C",x"0F",x"3C",x"0F",x"1E", -- 0x14F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1500
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1508
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1510
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1520
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1528
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1530
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1538
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1540
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1548
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1550
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1558
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1560
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1568
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1570
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1578
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1580
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1588
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1590
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1598
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15B8
		x"FF",x"FF",x"F1",x"F8",x"F7",x"F8",x"F0",x"F3", -- 0x15C0
		x"F0",x"F3",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x15C8
		x"F7",x"FE",x"F0",x"F0",x"FF",x"FF",x"F0",x"F0", -- 0x15D0
		x"F0",x"F0",x"F7",x"FE",x"F0",x"F0",x"FF",x"FF", -- 0x15D8
		x"FF",x"FF",x"F3",x"FF",x"F3",x"FF",x"FB",x"FF", -- 0x15E0
		x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x15F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1600
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1608
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1610
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1618
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1620
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1628
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1630
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1640
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1658
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1660
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1668
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1680
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"CF", -- 0x1688
		x"FF",x"CF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x1690
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1698
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16A0
		x"FF",x"FF",x"7F",x"FF",x"7F",x"FF",x"3F",x"FF", -- 0x16A8
		x"1F",x"FF",x"3F",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x16B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x16C0
		x"FF",x"CF",x"FF",x"9E",x"FF",x"BC",x"FF",x"3C", -- 0x16C8
		x"FF",x"78",x"FF",x"3C",x"FF",x"9E",x"FF",x"CF", -- 0x16D0
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x16E0
		x"1F",x"FF",x"C3",x"FF",x"E1",x"FF",x"F0",x"7F", -- 0x16E8
		x"F0",x"7F",x"E1",x"7F",x"C3",x"FF",x"97",x"FF", -- 0x16F0
		x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x16F8
		x"FF",x"FF",x"FF",x"EF",x"FF",x"DF",x"FF",x"FF", -- 0x1700
		x"DF",x"6F",x"FF",x"9E",x"EF",x"BC",x"FF",x"3C", -- 0x1708
		x"FF",x"3C",x"FF",x"78",x"EF",x"BC",x"FF",x"9E", -- 0x1710
		x"EF",x"4F",x"FF",x"EF",x"FF",x"5F",x"FF",x"EF", -- 0x1718
		x"FF",x"FF",x"FF",x"7F",x"DF",x"FF",x"7F",x"FF", -- 0x1720
		x"1F",x"7F",x"E1",x"FF",x"F0",x"5F",x"F0",x"7F", -- 0x1728
		x"F0",x"3F",x"F0",x"2F",x"F0",x"3F",x"E1",x"7F", -- 0x1730
		x"C3",x"FF",x"1F",x"7F",x"7F",x"BF",x"FF",x"FF", -- 0x1738
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF", -- 0x1740
		x"FF",x"FF",x"FF",x"4F",x"FF",x"DE",x"FF",x"BE", -- 0x1748
		x"FF",x"7C",x"DF",x"9E",x"FF",x"FE",x"FF",x"DF", -- 0x1750
		x"FF",x"FF",x"FF",x"7F",x"FF",x"EF",x"FF",x"BF", -- 0x1758
		x"FF",x"FF",x"DF",x"FF",x"7F",x"7F",x"BF",x"FF", -- 0x1760
		x"5F",x"FF",x"EB",x"FF",x"D3",x"7F",x"E1",x"BF", -- 0x1768
		x"F1",x"7F",x"E1",x"FF",x"F1",x"7F",x"5F",x"FF", -- 0x1770
		x"BF",x"FF",x"7F",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x1778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1788
		x"FF",x"FF",x"FF",x"FF",x"F1",x"F8",x"F7",x"F8", -- 0x1790
		x"F7",x"FB",x"F0",x"F3",x"F0",x"F3",x"FF",x"FF", -- 0x1798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17A8
		x"FF",x"FF",x"FF",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x17B0
		x"FB",x"FF",x"FB",x"FF",x"FB",x"FF",x"FF",x"FF", -- 0x17B8
		x"F0",x"F0",x"F0",x"F0",x"F7",x"FE",x"F0",x"F0", -- 0x17C0
		x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"F7",x"FE", -- 0x17C8
		x"F0",x"F0",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x17D0
		x"F7",x"FE",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x17D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x17F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x1800
		x"AD",x"FF",x"F8",x"FF",x"78",x"FF",x"5A",x"FF", -- 0x1808
		x"0F",x"FF",x"78",x"B7",x"F8",x"F3",x"EF",x"B7", -- 0x1810
		x"7F",x"FF",x"3F",x"FF",x"96",x"D3",x"B7",x"F8", -- 0x1818
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1820
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1828
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1830
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1838
		x"DE",x"D3",x"FF",x"FF",x"7F",x"FF",x"7F",x"B7", -- 0x1840
		x"FC",x"F3",x"BC",x"B7",x"0F",x"FF",x"3C",x"FF", -- 0x1848
		x"3C",x"FF",x"BC",x"FF",x"AD",x"FF",x"DF",x"FF", -- 0x1850
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1858
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1860
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1868
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1870
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1878
		x"FF",x"FF",x"DF",x"FF",x"AD",x"FF",x"F8",x"FF", -- 0x1880
		x"5A",x"FF",x"0F",x"FF",x"0F",x"3F",x"F0",x"B7", -- 0x1888
		x"EF",x"3F",x"1F",x"FF",x"C3",x"7F",x"E1",x"3F", -- 0x1890
		x"F0",x"3F",x"F0",x"97",x"F0",x"97",x"F0",x"A7", -- 0x1898
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"FF", -- 0x18B8
		x"F0",x"4E",x"F0",x"2F",x"F0",x"97",x"87",x"B7", -- 0x18C0
		x"3F",x"3F",x"4F",x"7F",x"8F",x"FF",x"F8",x"B7", -- 0x18C8
		x"F0",x"F3",x"78",x"B7",x"0F",x"FF",x"3C",x"FF", -- 0x18D0
		x"BC",x"FF",x"AD",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x18D8
		x"61",x"7F",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x18F8
		x"FF",x"FF",x"DF",x"FF",x"AD",x"FF",x"F8",x"FF", -- 0x1900
		x"3C",x"FF",x"0F",x"FF",x"1F",x"FF",x"2F",x"7F", -- 0x1908
		x"AF",x"3D",x"FF",x"5B",x"FF",x"1F",x"FF",x"CF", -- 0x1910
		x"8F",x"CF",x"AD",x"6F",x"78",x"7F",x"78",x"6F", -- 0x1918
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1920
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1928
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1930
		x"FF",x"FF",x"FF",x"FF",x"DE",x"F3",x"8C",x"D3", -- 0x1938
		x"E1",x"5E",x"C3",x"DE",x"1F",x"EF",x"FF",x"BF", -- 0x1940
		x"5E",x"5B",x"0F",x"3F",x"B7",x"FF",x"B7",x"F9", -- 0x1948
		x"C7",x"79",x"FE",x"F7",x"DE",x"7F",x"CF",x"7F", -- 0x1950
		x"CF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1958
		x"0C",x"97",x"4F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x1960
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1968
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1978
		x"FB",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"EF", -- 0x1980
		x"FF",x"FF",x"DD",x"FF",x"6F",x"7F",x"7B",x"3F", -- 0x1988
		x"D3",x"FF",x"3F",x"BF",x"FF",x"5B",x"DD",x"1F", -- 0x1990
		x"DD",x"EE",x"2E",x"DD",x"5B",x"23",x"D3",x"CE", -- 0x1998
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x19A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x19A8
		x"CF",x"FF",x"FF",x"FF",x"77",x"FF",x"FF",x"FF", -- 0x19B0
		x"FF",x"FF",x"BB",x"FF",x"7F",x"3F",x"7F",x"5B", -- 0x19B8
		x"6E",x"DE",x"EE",x"EF",x"DD",x"67",x"33",x"98", -- 0x19C0
		x"6F",x"DE",x"5E",x"1F",x"6F",x"3B",x"BF",x"CC", -- 0x19C8
		x"7B",x"77",x"2E",x"DD",x"DD",x"76",x"77",x"DE", -- 0x19D0
		x"FF",x"9F",x"EF",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x19D8
		x"FF",x"BF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19E0
		x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7", -- 0x19E8
		x"EF",x"7F",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A28
		x"9F",x"FF",x"9F",x"2F",x"F0",x"3F",x"99",x"FF", -- 0x1A30
		x"9B",x"CF",x"BF",x"3C",x"BF",x"78",x"EF",x"F0", -- 0x1A38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A58
		x"EF",x"F1",x"EF",x"E1",x"BF",x"78",x"BF",x"BC", -- 0x1A60
		x"F0",x"CF",x"99",x"FF",x"9B",x"FF",x"FF",x"FF", -- 0x1A68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"FF",x"FC", -- 0x1A88
		x"FF",x"BC",x"FF",x"CC",x"FF",x"CD",x"FF",x"FC", -- 0x1A90
		x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AA8
		x"F7",x"F3",x"FE",x"E1",x"EF",x"C3",x"CF",x"1E", -- 0x1AB0
		x"CF",x"F0",x"9E",x"F0",x"BC",x"F0",x"BC",x"F0", -- 0x1AB8
		x"FF",x"FF",x"FF",x"EF",x"FF",x"EF",x"FF",x"EF", -- 0x1AC0
		x"FF",x"FC",x"FF",x"EE",x"FF",x"EE",x"FF",x"FF", -- 0x1AC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AD8
		x"BC",x"F0",x"9E",x"F0",x"0F",x"78",x"4F",x"3C", -- 0x1AE0
		x"E1",x"3C",x"47",x"0F",x"7F",x"8F",x"FF",x"FF", -- 0x1AE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7", -- 0x1B00
		x"FF",x"7B",x"EF",x"3C",x"FF",x"3F",x"FF",x"BF", -- 0x1B08
		x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"CF",x"EF", -- 0x1B10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B20
		x"CF",x"FF",x"BC",x"7F",x"CF",x"FF",x"FF",x"8F", -- 0x1B28
		x"FF",x"3C",x"FF",x"0F",x"E7",x"5B",x"F3",x"3F", -- 0x1B30
		x"7F",x"FF",x"8F",x"FF",x"2D",x"7F",x"78",x"3F", -- 0x1B38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B40
		x"DE",x"F7",x"CF",x"7B",x"CF",x"7F",x"CF",x"FF", -- 0x1B48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B58
		x"F0",x"A7",x"78",x"2F",x"AD",x"7F",x"8F",x"9F", -- 0x1B60
		x"FF",x"8F",x"FD",x"BC",x"69",x"78",x"9F",x"78", -- 0x1B68
		x"FF",x"AF",x"FF",x"DE",x"FF",x"CF",x"FF",x"FF", -- 0x1B70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1B80
		x"FE",x"FF",x"DE",x"FF",x"DF",x"FF",x"DF",x"FF", -- 0x1B88
		x"FF",x"FF",x"FF",x"EE",x"FF",x"EE",x"FF",x"F7", -- 0x1B90
		x"EF",x"DD",x"FF",x"FF",x"FB",x"FF",x"7B",x"BB", -- 0x1B98
		x"FF",x"FF",x"FE",x"FF",x"FB",x"FF",x"7F",x"EE", -- 0x1BA0
		x"FF",x"DD",x"FF",x"77",x"DD",x"DD",x"BB",x"AB", -- 0x1BA8
		x"EF",x"6F",x"FF",x"3F",x"BB",x"DD",x"CC",x"AB", -- 0x1BB0
		x"77",x"DF",x"FF",x"FF",x"AD",x"DD",x"78",x"5D", -- 0x1BB8
		x"6F",x"AB",x"EF",x"D5",x"FF",x"5D",x"FF",x"AE", -- 0x1BC0
		x"FF",x"FF",x"DF",x"FF",x"DE",x"FF",x"EF",x"FF", -- 0x1BC8
		x"FF",x"FF",x"FF",x"DF",x"FF",x"DE",x"EF",x"EF", -- 0x1BD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1BD8
		x"F0",x"7F",x"69",x"FF",x"1F",x"AA",x"FF",x"67", -- 0x1BE0
		x"FF",x"47",x"00",x"DE",x"FF",x"67",x"17",x"FF", -- 0x1BE8
		x"DE",x"99",x"EF",x"7F",x"DD",x"AA",x"F7",x"77", -- 0x1BF0
		x"FF",x"BF",x"BF",x"8F",x"FF",x"CF",x"FF",x"FF", -- 0x1BF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C78
		x"FF",x"FF",x"FD",x"FF",x"FE",x"F7",x"FE",x"C3", -- 0x1C80
		x"FF",x"F0",x"FF",x"F0",x"FF",x"F8",x"FF",x"F8", -- 0x1C88
		x"FF",x"F8",x"FF",x"F0",x"FF",x"F0",x"FE",x"C3", -- 0x1C90
		x"FE",x"F7",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C98
		x"FB",x"FF",x"7B",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x1CA0
		x"F3",x"FF",x"F1",x"FF",x"F0",x"7F",x"F0",x"F3", -- 0x1CA8
		x"F0",x"7F",x"F1",x"FF",x"F3",x"FF",x"F3",x"FF", -- 0x1CB0
		x"F3",x"FF",x"7B",x"FF",x"FB",x"FF",x"FF",x"FF", -- 0x1CB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"CF", -- 0x1CC0
		x"1F",x"8F",x"1F",x"3F",x"E1",x"3E",x"E1",x"7A", -- 0x1CC8
		x"E1",x"3E",x"0F",x"1F",x"1F",x"0F",x"1F",x"8F", -- 0x1CD0
		x"1F",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"FF", -- 0x1CE0
		x"0F",x"3F",x"FF",x"9F",x"F4",x"CB",x"F4",x"E9", -- 0x1CE8
		x"F4",x"CB",x"BF",x"0F",x"0F",x"1F",x"0F",x"3F", -- 0x1CF0
		x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF8
		x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D00
		x"FF",x"3F",x"FF",x"9F",x"FF",x"FF",x"DF",x"FF", -- 0x1D08
		x"FF",x"FF",x"FF",x"7F",x"7F",x"FF",x"DD",x"FF", -- 0x1D10
		x"DD",x"EE",x"EE",x"DD",x"BF",x"33",x"7F",x"CE", -- 0x1D18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x1D20
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x1D28
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"DF",x"FF", -- 0x1D30
		x"EF",x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"FF", -- 0x1D38
		x"EE",x"FF",x"EE",x"FF",x"DD",x"77",x"33",x"99", -- 0x1D40
		x"FF",x"7F",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x1D48
		x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"BF",x"DF", -- 0x1D50
		x"FF",x"7F",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x1D58
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"BF", -- 0x1D60
		x"BF",x"FF",x"FF",x"FF",x"FE",x"FF",x"CF",x"FF", -- 0x1D68
		x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x1D80
		x"DF",x"FF",x"FF",x"BF",x"FF",x"DF",x"BF",x"FF", -- 0x1D88
		x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"FF",x"EF", -- 0x1D90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DA8
		x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DB0
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"DF",x"FF", -- 0x1DB8
		x"3F",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DC0
		x"FF",x"FF",x"FF",x"7F",x"EF",x"FF",x"7F",x"EF", -- 0x1DC8
		x"FF",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DD0
		x"FF",x"BF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DD8
		x"FF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE0
		x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE8
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E08
		x"FF",x"FF",x"EF",x"FF",x"EF",x"4F",x"DE",x"87", -- 0x1E10
		x"EE",x"4F",x"EF",x"6F",x"EF",x"6F",x"EF",x"6F", -- 0x1E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"9F",x"FF", -- 0x1E28
		x"9F",x"FF",x"1F",x"FF",x"0F",x"FF",x"E1",x"FF", -- 0x1E30
		x"1F",x"FF",x"1F",x"FF",x"78",x"7F",x"F6",x"B7", -- 0x1E38
		x"EF",x"6F",x"EF",x"4F",x"DE",x"87",x"EF",x"4F", -- 0x1E40
		x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E58
		x"0F",x"7F",x"1F",x"FF",x"69",x"FF",x"0F",x"FF", -- 0x1E60
		x"1F",x"FF",x"1F",x"FF",x"9F",x"FF",x"9F",x"FF", -- 0x1E68
		x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1ED8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1EF8
		x"FF",x"FF",x"FF",x"DF",x"FF",x"FF",x"FF",x"7F", -- 0x1F00
		x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F08
		x"DF",x"EF",x"BF",x"DF",x"FF",x"7F",x"FF",x"7F", -- 0x1F10
		x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"FF",x"FF", -- 0x1F18
		x"FF",x"DF",x"FF",x"7F",x"FF",x"FF",x"9F",x"FF", -- 0x1F20
		x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x1F28
		x"FF",x"7F",x"FF",x"FF",x"BB",x"DD",x"CC",x"BB", -- 0x1F30
		x"77",x"FF",x"FF",x"FF",x"FF",x"DD",x"DF",x"DD", -- 0x1F38
		x"FF",x"BB",x"FF",x"FF",x"BF",x"FF",x"BF",x"EE", -- 0x1F40
		x"DF",x"FF",x"FF",x"DF",x"FF",x"6F",x"FF",x"FF", -- 0x1F48
		x"FF",x"FF",x"FF",x"7F",x"FF",x"7F",x"FF",x"9F", -- 0x1F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F58
		x"9F",x"FF",x"FF",x"FF",x"FF",x"AA",x"FF",x"77", -- 0x1F60
		x"FF",x"77",x"CC",x"EF",x"FF",x"77",x"FF",x"FF", -- 0x1F68
		x"FF",x"FF",x"BF",x"FF",x"DF",x"FF",x"FF",x"DF", -- 0x1F70
		x"FF",x"FF",x"DF",x"FF",x"FF",x"9F",x"FF",x"FF", -- 0x1F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1F80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF", -- 0x1F88
		x"FF",x"FF",x"FF",x"DF",x"FF",x"BF",x"FF",x"FF", -- 0x1F90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF", -- 0x1F98
		x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"BF",x"DF", -- 0x1FA0
		x"FF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FA8
		x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FB0
		x"FF",x"EE",x"DF",x"FF",x"BF",x"FF",x"FF",x"FF", -- 0x1FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"7F", -- 0x1FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF", -- 0x1FC8
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD8
		x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF", -- 0x1FE0
		x"FF",x"FF",x"7F",x"FF",x"BF",x"DF",x"FF",x"FF", -- 0x1FE8
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x1FF0
		x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FF8
		x"FD",x"FF",x"D8",x"FF",x"88",x"FF",x"88",x"FF", -- 0x2000
		x"88",x"FF",x"80",x"FF",x"00",x"FF",x"00",x"DF", -- 0x2008
		x"00",x"DF",x"00",x"13",x"00",x"13",x"00",x"73", -- 0x2010
		x"00",x"FF",x"00",x"FF",x"00",x"10",x"11",x"CC", -- 0x2018
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2020
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2028
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2030
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"F3",x"FF", -- 0x2038
		x"F0",x"F0",x"00",x"DF",x"00",x"DF",x"00",x"13", -- 0x2040
		x"00",x"13",x"00",x"73",x"00",x"FF",x"00",x"FF", -- 0x2048
		x"00",x"FF",x"80",x"FF",x"88",x"FF",x"88",x"FF", -- 0x2050
		x"88",x"FF",x"D8",x"FF",x"FD",x"FF",x"FF",x"FF", -- 0x2058
		x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2060
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2068
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2070
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2078
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2080
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2088
		x"FF",x"FF",x"FF",x"FB",x"FF",x"B1",x"FF",x"11", -- 0x2090
		x"FF",x"11",x"FF",x"10",x"FF",x"00",x"EE",x"00", -- 0x2098
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20A8
		x"FF",x"FF",x"FF",x"FE",x"FF",x"EC",x"FF",x"EE", -- 0x20B0
		x"FF",x"EE",x"FF",x"EC",x"E8",x"00",x"00",x"33", -- 0x20B8
		x"FF",x"00",x"FF",x"10",x"FF",x"11",x"FF",x"11", -- 0x20C0
		x"FF",x"B1",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF", -- 0x20C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20D8
		x"F8",x"F0",x"FF",x"CC",x"FF",x"EE",x"FF",x"EE", -- 0x20E0
		x"FF",x"EC",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF", -- 0x20E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x20F8
		x"FF",x"FF",x"F7",x"FF",x"F7",x"FF",x"77",x"FF", -- 0x2100
		x"73",x"FF",x"63",x"FF",x"33",x"7F",x"30",x"BF", -- 0x2108
		x"40",x"F7",x"80",x"F7",x"20",x"FF",x"80",x"F8", -- 0x2110
		x"10",x"80",x"60",x"DC",x"91",x"70",x"00",x"A3", -- 0x2118
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2120
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2128
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x2130
		x"F7",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2138
		x"20",x"F3",x"A0",x"50",x"C0",x"80",x"E8",x"10", -- 0x2140
		x"C8",x"51",x"70",x"31",x"FC",x"11",x"FE",x"10", -- 0x2148
		x"FE",x"90",x"FF",x"90",x"FF",x"C8",x"FF",x"EC", -- 0x2150
		x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2158
		x"7F",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2160
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2168
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x2170
		x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2178
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2180
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2188
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2190
		x"FF",x"FF",x"FF",x"FF",x"FE",x"F7",x"EE",x"73", -- 0x2198
		x"FF",x"FE",x"FF",x"EC",x"FF",x"EC",x"FF",x"EC", -- 0x21A0
		x"FF",x"EC",x"FF",x"EC",x"FF",x"EC",x"FF",x"EC", -- 0x21A8
		x"FF",x"FE",x"FF",x"FE",x"FF",x"F8",x"FF",x"B8", -- 0x21B0
		x"FF",x"FE",x"FF",x"EC",x"FF",x"FC",x"FF",x"E8", -- 0x21B8
		x"FE",x"31",x"FE",x"10",x"FF",x"10",x"FF",x"80", -- 0x21C0
		x"FF",x"88",x"FF",x"10",x"FF",x"88",x"FF",x"CC", -- 0x21C8
		x"FF",x"EC",x"FF",x"FE",x"FF",x"FE",x"FF",x"FF", -- 0x21D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x21D8
		x"FF",x"D1",x"FC",x"00",x"D0",x"C0",x"F0",x"FF", -- 0x21E0
		x"F7",x"FF",x"F7",x"FF",x"F7",x"FF",x"73",x"FF", -- 0x21E8
		x"73",x"FF",x"73",x"FF",x"F3",x"FF",x"FF",x"FF", -- 0x21F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x21F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x2200
		x"BF",x"FF",x"D7",x"FF",x"F3",x"FF",x"71",x"FF", -- 0x2208
		x"F3",x"F1",x"F6",x"91",x"70",x"31",x"60",x"31", -- 0x2210
		x"D1",x"63",x"A2",x"77",x"44",x"F6",x"10",x"60", -- 0x2218
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2220
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2228
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2230
		x"FF",x"FF",x"7F",x"FF",x"37",x"FF",x"73",x"FF", -- 0x2238
		x"60",x"40",x"C0",x"80",x"90",x"00",x"F6",x"80", -- 0x2240
		x"FF",x"00",x"FE",x"FC",x"FF",x"FF",x"FF",x"FF", -- 0x2248
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2250
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2258
		x"73",x"FF",x"F7",x"FF",x"77",x"FF",x"73",x"FF", -- 0x2260
		x"31",x"FF",x"10",x"FF",x"D0",x"FF",x"FC",x"FF", -- 0x2268
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2270
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2278
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2280
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2288
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2290
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2298
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F3",x"FF", -- 0x22A0
		x"B1",x"FF",x"C0",x"FF",x"C8",x"76",x"E8",x"30", -- 0x22A8
		x"EC",x"00",x"FC",x"40",x"FE",x"80",x"FE",x"00", -- 0x22B0
		x"FE",x"40",x"FE",x"90",x"FF",x"F8",x"FF",x"E8", -- 0x22B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22C0
		x"FF",x"F9",x"FF",x"B0",x"FF",x"C0",x"FF",x"C8", -- 0x22C8
		x"FF",x"EC",x"FF",x"FE",x"FF",x"DD",x"FF",x"FF", -- 0x22D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22D8
		x"FF",x"D9",x"FF",x"EA",x"FF",x"98",x"FF",x"B0", -- 0x22E0
		x"FE",x"73",x"E4",x"F7",x"50",x"FF",x"31",x"FF", -- 0x22E8
		x"50",x"FF",x"90",x"FF",x"80",x"F7",x"C8",x"F7", -- 0x22F0
		x"FC",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x22F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2300
		x"FF",x"FF",x"FF",x"FF",x"FC",x"F7",x"E8",x"F7", -- 0x2308
		x"C8",x"F7",x"F2",x"F7",x"B2",x"FF",x"D4",x"BF", -- 0x2310
		x"10",x"DF",x"20",x"E5",x"40",x"40",x"40",x"80", -- 0x2318
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2320
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2328
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2330
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2338
		x"80",x"80",x"90",x"00",x"F0",x"00",x"EE",x"F0", -- 0x2340
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2348
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2350
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2358
		x"F3",x"FF",x"30",x"FF",x"10",x"F7",x"80",x"F7", -- 0x2360
		x"F8",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2368
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2370
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2378
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2380
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"D8", -- 0x2388
		x"FF",x"E8",x"FF",x"EC",x"FF",x"FC",x"FF",x"FE", -- 0x2390
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2398
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"F7",x"9F", -- 0x23A8
		x"31",x"F1",x"00",x"91",x"00",x"90",x"90",x"10", -- 0x23B0
		x"D0",x"10",x"F8",x"30",x"FC",x"20",x"EE",x"A0", -- 0x23B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"FF",x"EC", -- 0x23C8
		x"FF",x"EC",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x23D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23D8
		x"FF",x"D9",x"FF",x"C8",x"FF",x"88",x"FF",x"91", -- 0x23E0
		x"FF",x"B1",x"FF",x"33",x"F0",x"73",x"20",x"77", -- 0x23E8
		x"20",x"F3",x"C0",x"F1",x"C0",x"31",x"E8",x"10", -- 0x23F0
		x"BB",x"B0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x23F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2400
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FF", -- 0x2408
		x"F7",x"FF",x"47",x"7F",x"76",x"73",x"76",x"33", -- 0x2410
		x"10",x"00",x"10",x"00",x"10",x"00",x"00",x"00", -- 0x2418
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2420
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2428
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2430
		x"31",x"FF",x"10",x"FF",x"31",x"FF",x"F7",x"FF", -- 0x2438
		x"00",x"73",x"73",x"F7",x"77",x"FF",x"77",x"FF", -- 0x2440
		x"F7",x"FF",x"F7",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x2448
		x"FF",x"FF",x"FF",x"FF",x"73",x"FF",x"10",x"FF", -- 0x2450
		x"00",x"F7",x"10",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2458
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2460
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2468
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2470
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2478
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2480
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2488
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2490
		x"FF",x"80",x"FE",x"00",x"FF",x"80",x"FF",x"EC", -- 0x2498
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FC", -- 0x24A8
		x"FF",x"EC",x"1F",x"EC",x"C8",x"FD",x"C8",x"FD", -- 0x24B0
		x"40",x"31",x"40",x"20",x"40",x"20",x"80",x"20", -- 0x24B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x24D8
		x"88",x"31",x"FD",x"B9",x"FF",x"EC",x"FF",x"EC", -- 0x24E0
		x"FF",x"EC",x"FF",x"EC",x"FF",x"EC",x"FF",x"CC", -- 0x24E8
		x"FF",x"EE",x"FF",x"EE",x"FF",x"C8",x"FE",x"00", -- 0x24F0
		x"EC",x"00",x"FE",x"00",x"FF",x"EE",x"FF",x"FF", -- 0x24F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2500
		x"FF",x"FF",x"7B",x"FC",x"F1",x"C0",x"B0",x"00", -- 0x2508
		x"80",x"10",x"40",x"10",x"C0",x"31",x"20",x"F1", -- 0x2510
		x"70",x"F3",x"90",x"F7",x"00",x"77",x"71",x"FF", -- 0x2518
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2520
		x"FF",x"FF",x"F7",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x2528
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2530
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2538
		x"FB",x"FF",x"F3",x"FF",x"B1",x"FF",x"B1",x"FF", -- 0x2540
		x"D9",x"FF",x"D8",x"FF",x"FC",x"FC",x"EC",x"00", -- 0x2548
		x"EE",x"00",x"C8",x"30",x"80",x"71",x"20",x"33", -- 0x2550
		x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2558
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2560
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"77",x"FF", -- 0x2568
		x"F7",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2570
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2578
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2580
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2588
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"CF", -- 0x2590
		x"FF",x"BE",x"FF",x"FE",x"FF",x"FF",x"FF",x"FE", -- 0x2598
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25A0
		x"FF",x"FF",x"FF",x"EF",x"EC",x"D7",x"EC",x"73", -- 0x25A8
		x"DC",x"31",x"FE",x"31",x"EE",x"D4",x"72",x"C0", -- 0x25B0
		x"20",x"62",x"00",x"60",x"90",x"20",x"40",x"30", -- 0x25B8
		x"FF",x"EC",x"FF",x"C8",x"FF",x"80",x"FE",x"00", -- 0x25C0
		x"EE",x"30",x"FE",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x25C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25D8
		x"60",x"90",x"30",x"10",x"10",x"E0",x"71",x"77", -- 0x25E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x25F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"71", -- 0x2600
		x"EE",x"31",x"CC",x"73",x"88",x"73",x"80",x"77", -- 0x2608
		x"00",x"F7",x"00",x"F7",x"90",x"FF",x"50",x"FF", -- 0x2610
		x"00",x"FF",x"30",x"FF",x"73",x"FF",x"73",x"FF", -- 0x2618
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2620
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2628
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2630
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2638
		x"B9",x"FF",x"91",x"FF",x"20",x"FF",x"FE",x"74", -- 0x2640
		x"FF",x"80",x"FF",x"80",x"FF",x"80",x"FF",x"C0", -- 0x2648
		x"FF",x"A0",x"FF",x"B1",x"FF",x"B3",x"FF",x"F7", -- 0x2650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2658
		x"FF",x"FF",x"FF",x"FF",x"F1",x"FF",x"31",x"FF", -- 0x2660
		x"31",x"FF",x"33",x"FF",x"77",x"FF",x"77",x"FF", -- 0x2668
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2670
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2678
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2680
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2688
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2690
		x"FF",x"FF",x"FF",x"CF",x"FF",x"BF",x"FF",x"FE", -- 0x2698
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"1D",x"EF",x"C8", -- 0x26A8
		x"F1",x"E8",x"90",x"DC",x"C0",x"50",x"F9",x"00", -- 0x26B0
		x"EC",x"88",x"D4",x"44",x"40",x"80",x"20",x"51", -- 0x26B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"EE", -- 0x26C0
		x"FF",x"CC",x"FF",x"C8",x"FF",x"80",x"FF",x"F0", -- 0x26C8
		x"FF",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26D8
		x"80",x"20",x"40",x"C0",x"20",x"70",x"00",x"B3", -- 0x26E0
		x"10",x"F7",x"33",x"FF",x"F7",x"FF",x"FF",x"FF", -- 0x26E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x26F8
		x"FF",x"FF",x"F9",x"FF",x"91",x"FF",x"B1",x"FF", -- 0x2700
		x"31",x"FF",x"31",x"FF",x"31",x"FF",x"31",x"FF", -- 0x2708
		x"33",x"FF",x"73",x"FF",x"73",x"FF",x"73",x"FF", -- 0x2710
		x"51",x"FF",x"33",x"FF",x"33",x"FF",x"71",x"FF", -- 0x2718
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2720
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2728
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2730
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2738
		x"B8",x"FF",x"90",x"F7",x"F0",x"71",x"FE",x"80", -- 0x2740
		x"FF",x"CC",x"FF",x"EE",x"FF",x"EC",x"FF",x"EC", -- 0x2748
		x"FF",x"CC",x"FF",x"CC",x"FF",x"CC",x"FF",x"FF", -- 0x2750
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2758
		x"C8",x"FF",x"C8",x"FF",x"80",x"FF",x"10",x"FF", -- 0x2760
		x"11",x"FF",x"11",x"FF",x"20",x"FF",x"B3",x"FF", -- 0x2768
		x"73",x"FF",x"77",x"FF",x"F7",x"FF",x"FF",x"FF", -- 0x2770
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2778
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2788
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EC", -- 0x2790
		x"FF",x"CC",x"FF",x"EC",x"FF",x"FE",x"FF",x"FF", -- 0x2798
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27A0
		x"FF",x"FE",x"FF",x"FE",x"DE",x"F4",x"CE",x"60", -- 0x27A8
		x"BC",x"20",x"FE",x"90",x"FF",x"40",x"F3",x"90", -- 0x27B0
		x"30",x"00",x"66",x"00",x"D1",x"00",x"F8",x"80", -- 0x27B8
		x"FF",x"FF",x"FF",x"FE",x"FF",x"CE",x"FF",x"CE", -- 0x27C0
		x"FF",x"BC",x"FF",x"EE",x"FF",x"FF",x"FF",x"FE", -- 0x27C8
		x"FF",x"EE",x"FF",x"EC",x"FF",x"FC",x"FF",x"FF", -- 0x27D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27D8
		x"CC",x"E0",x"D8",x"30",x"C0",x"40",x"20",x"30", -- 0x27E0
		x"10",x"31",x"60",x"F3",x"10",x"B3",x"00",x"FF", -- 0x27E8
		x"31",x"FF",x"F3",x"FF",x"F7",x"FF",x"FF",x"FF", -- 0x27F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x27F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2800
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2808
		x"FF",x"FF",x"F7",x"FF",x"73",x"FF",x"77",x"FF", -- 0x2810
		x"77",x"FF",x"73",x"FF",x"00",x"71",x"CC",x"00", -- 0x2818
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2820
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2828
		x"FF",x"FF",x"FD",x"FF",x"D8",x"FF",x"88",x"FF", -- 0x2830
		x"88",x"FF",x"80",x"FF",x"00",x"FF",x"00",x"77", -- 0x2838
		x"F0",x"F1",x"33",x"FF",x"77",x"FF",x"77",x"FF", -- 0x2840
		x"73",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2848
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2850
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2858
		x"00",x"FF",x"00",x"FF",x"88",x"FF",x"88",x"FF", -- 0x2860
		x"D8",x"FF",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2868
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2870
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2878
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2880
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2888
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2890
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FC", -- 0x2898
		x"FF",x"FB",x"FF",x"B1",x"FF",x"11",x"FF",x"11", -- 0x28A0
		x"FF",x"11",x"FF",x"10",x"FF",x"00",x"FF",x"00", -- 0x28A8
		x"FF",x"00",x"CC",x"00",x"8C",x"00",x"AC",x"00", -- 0x28B0
		x"BF",x"00",x"BF",x"00",x"80",x"00",x"33",x"88", -- 0x28B8
		x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x28D8
		x"F0",x"F0",x"FF",x"00",x"FF",x"00",x"CC",x"00", -- 0x28E0
		x"8C",x"00",x"AC",x"00",x"BF",x"00",x"BF",x"00", -- 0x28E8
		x"FF",x"00",x"FF",x"10",x"FF",x"11",x"FF",x"11", -- 0x28F0
		x"FF",x"11",x"FF",x"B1",x"FF",x"FB",x"FF",x"FF", -- 0x28F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2900
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FE", -- 0x2908
		x"FF",x"FE",x"FF",x"FE",x"FF",x"FE",x"FF",x"FC", -- 0x2910
		x"FF",x"C0",x"E8",x"20",x"C0",x"F3",x"B8",x"FF", -- 0x2918
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2920
		x"FF",x"FF",x"FF",x"FF",x"73",x"FF",x"73",x"FF", -- 0x2928
		x"31",x"FF",x"31",x"FF",x"00",x"FF",x"11",x"FF", -- 0x2930
		x"10",x"FF",x"80",x"F7",x"C0",x"F7",x"E8",x"77", -- 0x2938
		x"F1",x"FF",x"F7",x"FF",x"77",x"FF",x"F7",x"FF", -- 0x2940
		x"D1",x"FF",x"F1",x"FF",x"77",x"FF",x"F7",x"FF", -- 0x2948
		x"73",x"FF",x"73",x"FF",x"73",x"FF",x"73",x"FF", -- 0x2950
		x"73",x"FF",x"33",x"FF",x"73",x"FF",x"F3",x"FF", -- 0x2958
		x"FC",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2960
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2968
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2978
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x2980
		x"FF",x"FE",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x2988
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2990
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF", -- 0x2998
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FF", -- 0x29A0
		x"73",x"FF",x"31",x"FF",x"30",x"FF",x"90",x"FF", -- 0x29A8
		x"80",x"F7",x"80",x"F3",x"88",x"60",x"E8",x"11", -- 0x29B0
		x"80",x"51",x"10",x"10",x"80",x"10",x"4C",x"60", -- 0x29B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x29C0
		x"FF",x"EE",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x29C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x29D8
		x"BC",x"80",x"C8",x"98",x"B3",x"60",x"10",x"80", -- 0x29E0
		x"71",x"00",x"F3",x"20",x"FE",x"90",x"FF",x"00", -- 0x29E8
		x"EF",x"80",x"FF",x"4C",x"FF",x"AC",x"FF",x"EC", -- 0x29F0
		x"FF",x"EE",x"FF",x"FE",x"FF",x"FE",x"FF",x"FF", -- 0x29F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"73", -- 0x2A00
		x"FE",x"31",x"FE",x"30",x"FE",x"00",x"FF",x"80", -- 0x2A08
		x"FF",x"C0",x"FF",x"A0",x"FE",x"70",x"CC",x"F6", -- 0x2A10
		x"88",x"F7",x"90",x"FF",x"20",x"FF",x"F9",x"FF", -- 0x2A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A20
		x"FF",x"FF",x"77",x"FF",x"F7",x"FF",x"73",x"FF", -- 0x2A28
		x"71",x"FF",x"31",x"FF",x"31",x"FF",x"F1",x"FF", -- 0x2A30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A38
		x"71",x"FF",x"D1",x"FF",x"F1",x"FF",x"B1",x"77", -- 0x2A40
		x"70",x"FF",x"90",x"FF",x"30",x"F7",x"40",x"F7", -- 0x2A48
		x"C0",x"73",x"C0",x"73",x"EC",x"71",x"FE",x"31", -- 0x2A50
		x"FF",x"31",x"FF",x"F9",x"FF",x"FF",x"FF",x"FF", -- 0x2A58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2A88
		x"FF",x"B0",x"FF",x"C0",x"FF",x"C8",x"FF",x"E8", -- 0x2A90
		x"FF",x"FC",x"FF",x"FE",x"FF",x"FF",x"FF",x"FE", -- 0x2A98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AA8
		x"FF",x"FF",x"F3",x"FF",x"71",x"FF",x"30",x"BB", -- 0x2AB0
		x"00",x"F7",x"A0",x"F0",x"D0",x"90",x"B0",x"20", -- 0x2AB8
		x"FF",x"FE",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x2AC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AD8
		x"60",x"51",x"64",x"80",x"7E",x"10",x"AC",x"74", -- 0x2AE0
		x"C8",x"F8",x"D9",x"E0",x"98",x"F4",x"F8",x"FC", -- 0x2AE8
		x"FF",x"E8",x"FF",x"D8",x"FF",x"BD",x"FF",x"DF", -- 0x2AF0
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2AF8
		x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"88",x"D5", -- 0x2B00
		x"88",x"31",x"C8",x"90",x"EC",x"80",x"FC",x"00", -- 0x2B08
		x"EE",x"E0",x"EC",x"F0",x"CC",x"FF",x"D8",x"FF", -- 0x2B10
		x"98",x"FF",x"91",x"FF",x"31",x"FF",x"B9",x"FF", -- 0x2B18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B20
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"77",x"FF", -- 0x2B28
		x"77",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B38
		x"10",x"77",x"10",x"F7",x"10",x"F3",x"20",x"B1", -- 0x2B40
		x"C0",x"90",x"D8",x"00",x"D8",x"00",x"D8",x"C8", -- 0x2B48
		x"9F",x"FC",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B60
		x"FF",x"FF",x"F7",x"FF",x"73",x"FF",x"73",x"FF", -- 0x2B68
		x"33",x"FF",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2B90
		x"FE",x"10",x"FE",x"00",x"FE",x"80",x"FF",x"E0", -- 0x2B98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BB0
		x"F7",x"77",x"00",x"90",x"20",x"10",x"20",x"10", -- 0x2BB8
		x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BD8
		x"40",x"20",x"C0",x"20",x"90",x"51",x"B1",x"E2", -- 0x2BE0
		x"B1",x"EA",x"3F",x"90",x"DF",x"91",x"FF",x"B1", -- 0x2BE8
		x"FF",x"71",x"FF",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x2BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2BF8
		x"FF",x"FF",x"FF",x"FF",x"00",x"F7",x"00",x"73", -- 0x2C00
		x"00",x"F7",x"10",x"FF",x"F3",x"FF",x"FF",x"FF", -- 0x2C08
		x"F7",x"FF",x"F7",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x2C10
		x"77",x"FF",x"73",x"FF",x"31",x"77",x"00",x"71", -- 0x2C18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C38
		x"00",x"00",x"10",x"00",x"10",x"00",x"00",x"00", -- 0x2C40
		x"66",x"33",x"76",x"33",x"77",x"1F",x"F7",x"FF", -- 0x2C48
		x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C58
		x"73",x"FF",x"10",x"FF",x"00",x"F7",x"10",x"FF", -- 0x2C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2C98
		x"FF",x"FF",x"FF",x"EE",x"EC",x"00",x"C8",x"00", -- 0x2CA0
		x"EC",x"00",x"FE",x"00",x"FF",x"88",x"FF",x"EE", -- 0x2CA8
		x"FF",x"CC",x"FF",x"EC",x"FF",x"EC",x"FF",x"EC", -- 0x2CB0
		x"FF",x"EC",x"FF",x"A8",x"FD",x"31",x"80",x"B1", -- 0x2CB8
		x"FF",x"C8",x"FE",x"00",x"EC",x"00",x"FE",x"00", -- 0x2CC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CD8
		x"80",x"A0",x"00",x"20",x"00",x"20",x"00",x"31", -- 0x2CE0
		x"88",x"FD",x"C8",x"FD",x"CF",x"6C",x"FF",x"EC", -- 0x2CE8
		x"FF",x"FC",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x2CF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2CF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D10
		x"FF",x"FF",x"EE",x"E0",x"E0",x"00",x"60",x"00", -- 0x2D18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D30
		x"F8",x"FF",x"00",x"FF",x"10",x"FF",x"30",x"FF", -- 0x2D38
		x"10",x"00",x"00",x"10",x"00",x"90",x"00",x"C0", -- 0x2D40
		x"D4",x"D8",x"D4",x"EF",x"E2",x"FF",x"40",x"F7", -- 0x2D48
		x"68",x"F7",x"FC",x"F7",x"FE",x"F7",x"FF",x"FF", -- 0x2D50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D58
		x"F3",x"FF",x"F7",x"FF",x"FF",x"FF",x"BF",x"FF", -- 0x2D60
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D80
		x"FF",x"FF",x"FF",x"EC",x"FF",x"C8",x"FF",x"80", -- 0x2D88
		x"FF",x"80",x"FF",x"F1",x"FF",x"FF",x"FF",x"FF", -- 0x2D90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2D98
		x"FF",x"FF",x"FF",x"F1",x"FE",x"31",x"44",x"71", -- 0x2DA0
		x"00",x"73",x"00",x"F3",x"00",x"F7",x"10",x"FF", -- 0x2DA8
		x"E4",x"FF",x"EC",x"F7",x"FE",x"73",x"FE",x"33", -- 0x2DB0
		x"FF",x"B1",x"FF",x"90",x"FF",x"40",x"FF",x"40", -- 0x2DB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DC0
		x"FF",x"FF",x"FF",x"FE",x"FF",x"EC",x"FF",x"C8", -- 0x2DC8
		x"FF",x"C8",x"FF",x"D8",x"FF",x"FF",x"FF",x"FF", -- 0x2DD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DD8
		x"FF",x"B1",x"BA",x"A0",x"F8",x"10",x"88",x"90", -- 0x2DE0
		x"E0",x"80",x"20",x"40",x"10",x"31",x"10",x"31", -- 0x2DE8
		x"60",x"B1",x"F7",x"E1",x"FF",x"DF",x"FF",x"FF", -- 0x2DF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE", -- 0x2E08
		x"FF",x"EC",x"FF",x"C0",x"B8",x"80",x"A8",x"00", -- 0x2E10
		x"C0",x"10",x"90",x"10",x"40",x"B1",x"20",x"50", -- 0x2E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E20
		x"FF",x"FF",x"FF",x"FF",x"F1",x"FF",x"31",x"FF", -- 0x2E28
		x"71",x"FF",x"73",x"FF",x"F3",x"FF",x"F7",x"FF", -- 0x2E30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x2E38
		x"98",x"60",x"00",x"F5",x"A2",x"F7",x"51",x"33", -- 0x2E40
		x"20",x"31",x"72",x"31",x"23",x"91",x"D3",x"F9", -- 0x2E48
		x"37",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E58
		x"BF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E80
		x"FF",x"DC",x"FF",x"EE",x"FF",x"CC",x"FF",x"88", -- 0x2E88
		x"FF",x"80",x"FF",x"90",x"FE",x"30",x"FE",x"F3", -- 0x2E90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2E98
		x"FF",x"FF",x"FC",x"F7",x"D8",x"F7",x"80",x"FF", -- 0x2EA0
		x"10",x"FF",x"10",x"FF",x"70",x"FF",x"11",x"FF", -- 0x2EA8
		x"91",x"FF",x"C0",x"F7",x"EC",x"73",x"FE",x"31", -- 0x2EB0
		x"FE",x"10",x"FF",x"80",x"FF",x"40",x"FF",x"A8", -- 0x2EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2ED8
		x"FF",x"98",x"EE",x"98",x"FF",x"C0",x"FF",x"00", -- 0x2EE0
		x"FE",x"00",x"FE",x"20",x"EC",x"10",x"EC",x"00", -- 0x2EE8
		x"C8",x"33",x"C8",x"77",x"C0",x"FF",x"91",x"FF", -- 0x2EF0
		x"F3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2EF8
		x"FF",x"FF",x"FF",x"F9",x"FF",x"F1",x"FF",x"91", -- 0x2F00
		x"FE",x"31",x"FE",x"31",x"EC",x"31",x"EC",x"33", -- 0x2F08
		x"C8",x"73",x"C0",x"71",x"80",x"10",x"10",x"01", -- 0x2F10
		x"30",x"61",x"00",x"F7",x"00",x"F3",x"00",x"71", -- 0x2F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F28
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x2F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F38
		x"11",x"98",x"40",x"44",x"50",x"80",x"11",x"F0", -- 0x2F40
		x"10",x"DF",x"00",x"B7",x"00",x"37",x"30",x"F7", -- 0x2F48
		x"33",x"FF",x"73",x"FF",x"73",x"FF",x"77",x"FF", -- 0x2F50
		x"77",x"FF",x"F7",x"FF",x"F7",x"FF",x"FF",x"FF", -- 0x2F58
		x"F7",x"FF",x"F3",x"FF",x"73",x"FF",x"F3",x"FF", -- 0x2F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2F80
		x"FF",x"FD",x"FF",x"D8",x"FF",x"98",x"FF",x"80", -- 0x2F88
		x"FF",x"80",x"EE",x"00",x"FF",x"00",x"FE",x"00", -- 0x2F90
		x"FE",x"00",x"FE",x"10",x"EE",x"31",x"FE",x"31", -- 0x2F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FA8
		x"FF",x"FF",x"FF",x"EE",x"FF",x"FF",x"F3",x"FE", -- 0x2FB0
		x"10",x"F4",x"E0",x"00",x"FC",x"22",x"FF",x"C0", -- 0x2FB8
		x"FE",x"73",x"FF",x"F3",x"FF",x"FF",x"FF",x"FF", -- 0x2FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x2FD8
		x"FF",x"D8",x"FF",x"DC",x"FF",x"CC",x"FF",x"CC", -- 0x2FE0
		x"FF",x"88",x"FF",x"FC",x"FF",x"CC",x"FF",x"CC", -- 0x2FE8
		x"FF",x"CC",x"FF",x"CC",x"FF",x"CC",x"FF",x"CC", -- 0x2FF0
		x"FF",x"CC",x"FF",x"CC",x"FF",x"EC",x"FF",x"FC", -- 0x2FF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3000
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3008
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3010
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3018
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3020
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3028
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3030
		x"FF",x"FF",x"FF",x"F8",x"FF",x"FE",x"FF",x"EF", -- 0x3038
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3040
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3048
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"F0",x"F0", -- 0x3050
		x"F0",x"F0",x"00",x"00",x"00",x"01",x"00",x"70", -- 0x3058
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3060
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3068
		x"FD",x"FF",x"FD",x"FF",x"69",x"F0",x"F0",x"F0", -- 0x3070
		x"F0",x"F0",x"00",x"00",x"84",x"00",x"C0",x"00", -- 0x3078
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3080
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3088
		x"FF",x"FF",x"FF",x"F8",x"FF",x"C0",x"FF",x"C0", -- 0x3090
		x"FE",x"C0",x"FE",x"C0",x"FE",x"C0",x"FE",x"C0", -- 0x3098
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x30A8
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"77",x"FF", -- 0x30B0
		x"73",x"FF",x"33",x"FF",x"33",x"FF",x"31",x"FF", -- 0x30B8
		x"FE",x"C0",x"FE",x"C0",x"FE",x"C0",x"FE",x"C0", -- 0x30C0
		x"FE",x"C0",x"FE",x"C0",x"FE",x"C0",x"FE",x"C0", -- 0x30C8
		x"FE",x"C0",x"FE",x"C0",x"FE",x"C0",x"FE",x"C0", -- 0x30D0
		x"3C",x"C0",x"68",x"C0",x"F0",x"00",x"3C",x"00", -- 0x30D8
		x"31",x"FF",x"31",x"FF",x"31",x"FF",x"30",x"FF", -- 0x30E0
		x"30",x"FF",x"30",x"FF",x"30",x"FF",x"30",x"FF", -- 0x30E8
		x"30",x"F7",x"30",x"F7",x"30",x"F7",x"30",x"F0", -- 0x30F0
		x"30",x"F0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3100
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3108
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3110
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3118
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3120
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3128
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3130
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3138
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3140
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3148
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3150
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3158
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3160
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3168
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3170
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3178
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3180
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3188
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3190
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3198
		x"FF",x"FE",x"FF",x"FE",x"FF",x"FE",x"FF",x"FE", -- 0x31A0
		x"FF",x"FE",x"FF",x"FE",x"FF",x"FC",x"FF",x"FC", -- 0x31A8
		x"FF",x"FC",x"FF",x"FC",x"FF",x"FC",x"FF",x"F8", -- 0x31B0
		x"FF",x"F8",x"FF",x"F8",x"FF",x"F8",x"FF",x"F0", -- 0x31B8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x31C8
		x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x31D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D8
		x"FF",x"F0",x"FF",x"F0",x"FF",x"F0",x"FE",x"F0", -- 0x31E0
		x"FE",x"F0",x"FE",x"F0",x"FC",x"F0",x"FC",x"F0", -- 0x31E8
		x"F8",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x31F0
		x"00",x"00",x"00",x"00",x"00",x"25",x"10",x"F0", -- 0x31F8
		x"FF",x"E0",x"FF",x"E0",x"FF",x"E0",x"FF",x"E0", -- 0x3200
		x"FE",x"E0",x"FE",x"E0",x"FE",x"E0",x"FE",x"E0", -- 0x3208
		x"FE",x"E0",x"FE",x"E0",x"FC",x"E0",x"FC",x"E0", -- 0x3210
		x"FC",x"E0",x"FC",x"E0",x"FC",x"E0",x"FC",x"E0", -- 0x3218
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3220
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3228
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3230
		x"00",x"30",x"00",x"30",x"00",x"C0",x"E0",x"00", -- 0x3238
		x"FC",x"E0",x"F8",x"E0",x"F8",x"E0",x"F8",x"E0", -- 0x3240
		x"F8",x"E0",x"F8",x"E0",x"F8",x"E0",x"F8",x"E0", -- 0x3248
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3250
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3258
		x"00",x"C0",x"F0",x"30",x"00",x"D0",x"00",x"60", -- 0x3260
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3268
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3270
		x"00",x"30",x"00",x"C0",x"E0",x"00",x"00",x"80", -- 0x3278
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3280
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3288
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3290
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3298
		x"F0",x"30",x"00",x"D0",x"00",x"60",x"00",x"30", -- 0x32A0
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x32A8
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x32B0
		x"00",x"40",x"70",x"00",x"00",x"40",x"70",x"90", -- 0x32B8
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x32C0
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x32C8
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x32D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D8
		x"00",x"E0",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x32E0
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x32E8
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x32F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10", -- 0x32F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3300
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3308
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3310
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3318
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3320
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3328
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F3", -- 0x3330
		x"FE",x"31",x"EC",x"31",x"CC",x"31",x"C8",x"31", -- 0x3338
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3340
		x"FF",x"FE",x"FF",x"EE",x"FF",x"EE",x"FF",x"EC", -- 0x3348
		x"FF",x"EC",x"FF",x"EC",x"FF",x"E8",x"FF",x"E8", -- 0x3350
		x"FF",x"E8",x"FF",x"E8",x"FF",x"E8",x"FF",x"E0", -- 0x3358
		x"88",x"31",x"80",x"31",x"00",x"31",x"00",x"31", -- 0x3360
		x"00",x"31",x"00",x"31",x"00",x"31",x"00",x"31", -- 0x3368
		x"00",x"31",x"00",x"31",x"00",x"31",x"00",x"31", -- 0x3370
		x"00",x"31",x"00",x"31",x"00",x"30",x"00",x"30", -- 0x3378
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3380
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3388
		x"FF",x"FF",x"F7",x"FF",x"F0",x"FF",x"F0",x"F3", -- 0x3390
		x"00",x"5A",x"00",x"10",x"80",x"A0",x"00",x"00", -- 0x3398
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33B0
		x"FF",x"FF",x"F7",x"FF",x"7F",x"FF",x"F7",x"FF", -- 0x33B8
		x"80",x"82",x"00",x"30",x"F0",x"5A",x"F0",x"F3", -- 0x33C0
		x"F0",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33D8
		x"7F",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x33F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3400
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3408
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3410
		x"F0",x"F3",x"F0",x"F1",x"00",x"10",x"00",x"10", -- 0x3418
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3420
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3428
		x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"BF",x"FF", -- 0x3430
		x"BF",x"FF",x"BF",x"FF",x"BF",x"FF",x"BF",x"FF", -- 0x3438
		x"00",x"10",x"F0",x"F0",x"F0",x"F1",x"F0",x"F3", -- 0x3440
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3448
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"F1", -- 0x3450
		x"F0",x"F0",x"00",x"10",x"00",x"00",x"00",x"00", -- 0x3458
		x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3460
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3468
		x"FF",x"FF",x"DF",x"FF",x"DF",x"FF",x"DF",x"FF", -- 0x3470
		x"DF",x"FF",x"D7",x"FF",x"D7",x"FF",x"87",x"FF", -- 0x3478
		x"F0",x"F0",x"F0",x"F0",x"F0",x"F1",x"FF",x"FF", -- 0x3480
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x3488
		x"F7",x"FF",x"F7",x"FF",x"F0",x"F0",x"F0",x"F0", -- 0x3490
		x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0", -- 0x3498
		x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34A8
		x"EF",x"FF",x"EF",x"FF",x"EF",x"FF",x"E7",x"FF", -- 0x34B0
		x"63",x"FF",x"63",x"FF",x"43",x"7F",x"F3",x"FF", -- 0x34B8
		x"F0",x"F0",x"70",x"F0",x"F7",x"FF",x"F7",x"FF", -- 0x34C0
		x"F7",x"FF",x"F7",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x34C8
		x"F7",x"FF",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x34D0
		x"00",x"00",x"00",x"00",x"25",x"00",x"F0",x"00", -- 0x34D8
		x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x34E8
		x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x34F0
		x"00",x"30",x"00",x"00",x"00",x"30",x"00",x"00", -- 0x34F8
		x"E0",x"00",x"84",x"00",x"08",x"00",x"EE",x"10", -- 0x3500
		x"EE",x"30",x"EE",x"60",x"EE",x"C0",x"FE",x"C0", -- 0x3508
		x"FE",x"C0",x"FE",x"C0",x"FE",x"C0",x"FE",x"C0", -- 0x3510
		x"FE",x"C0",x"FE",x"C0",x"FE",x"C0",x"FE",x"C0", -- 0x3518
		x"10",x"80",x"70",x"F0",x"F0",x"F0",x"B0",x"F0", -- 0x3520
		x"30",x"F7",x"30",x"F7",x"30",x"F7",x"30",x"FF", -- 0x3528
		x"30",x"FF",x"30",x"FF",x"30",x"FF",x"30",x"FF", -- 0x3530
		x"31",x"FF",x"31",x"FF",x"31",x"FF",x"31",x"FF", -- 0x3538
		x"FE",x"C0",x"FE",x"C0",x"FE",x"C0",x"FF",x"C0", -- 0x3540
		x"FF",x"C0",x"FF",x"F8",x"FF",x"FF",x"FF",x"FF", -- 0x3548
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3550
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3558
		x"33",x"FF",x"33",x"FF",x"73",x"FF",x"77",x"FF", -- 0x3560
		x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3568
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3570
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3578
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3580
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3588
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3590
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3598
		x"FF",x"FE",x"FF",x"F8",x"FF",x"FF",x"FF",x"FF", -- 0x35A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35B0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35B8
		x"00",x"01",x"F0",x"C0",x"F0",x"F0",x"F0",x"F0", -- 0x35C0
		x"FF",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35D8
		x"84",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x35E0
		x"0F",x"F0",x"BD",x"FF",x"FD",x"FF",x"FF",x"FF", -- 0x35E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x35F8
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x3600
		x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x3608
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3610
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3618
		x"00",x"25",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x3620
		x"F0",x"80",x"C0",x"00",x"88",x"30",x"CC",x"F0", -- 0x3628
		x"DC",x"F0",x"FE",x"F0",x"FE",x"F0",x"FE",x"F0", -- 0x3630
		x"FF",x"F0",x"FF",x"F0",x"FF",x"F0",x"FF",x"F0", -- 0x3638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3640
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3648
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3658
		x"FF",x"F8",x"FF",x"F8",x"FF",x"F8",x"FF",x"F8", -- 0x3660
		x"FF",x"FC",x"FF",x"FC",x"FF",x"FC",x"FF",x"FC", -- 0x3668
		x"FF",x"FC",x"FF",x"FE",x"FF",x"FE",x"FF",x"FE", -- 0x3670
		x"FF",x"FE",x"FF",x"FE",x"FF",x"FE",x"FF",x"FF", -- 0x3678
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3680
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3688
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3690
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3698
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F8
		x"00",x"00",x"00",x"00",x"F0",x"E0",x"E0",x"00", -- 0x3700
		x"00",x"70",x"70",x"F0",x"F0",x"F0",x"F0",x"E0", -- 0x3708
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3710
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3718
		x"00",x"00",x"00",x"00",x"00",x"F0",x"E0",x"00", -- 0x3720
		x"F0",x"E0",x"C0",x"70",x"00",x"30",x"00",x"30", -- 0x3728
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3730
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3738
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3740
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3748
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3750
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3758
		x"00",x"40",x"70",x"00",x"00",x"70",x"70",x"80", -- 0x3760
		x"00",x"70",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3768
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x3770
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"40", -- 0x3778
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F0",x"E0", -- 0x3780
		x"F0",x"E0",x"F0",x"E0",x"F0",x"E0",x"F8",x"E0", -- 0x3788
		x"F8",x"E0",x"F8",x"E0",x"F8",x"E0",x"F8",x"E0", -- 0x3790
		x"F8",x"E0",x"F8",x"E0",x"FC",x"E0",x"FC",x"E0", -- 0x3798
		x"E0",x"00",x"00",x"F0",x"F0",x"10",x"00",x"E0", -- 0x37A0
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x37A8
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x37B0
		x"00",x"30",x"00",x"20",x"00",x"80",x"E0",x"00", -- 0x37B8
		x"FC",x"E0",x"FC",x"E0",x"FC",x"E0",x"FC",x"E0", -- 0x37C0
		x"FC",x"E0",x"FE",x"E0",x"FE",x"E0",x"FE",x"E0", -- 0x37C8
		x"FE",x"E0",x"FE",x"E0",x"FE",x"E0",x"FF",x"E0", -- 0x37D0
		x"FF",x"E0",x"FF",x"E0",x"FF",x"E0",x"FF",x"E0", -- 0x37D8
		x"00",x"F0",x"F0",x"10",x"00",x"E0",x"00",x"30", -- 0x37E0
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x37E8
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x37F0
		x"00",x"30",x"00",x"30",x"00",x"30",x"00",x"30", -- 0x37F8
		x"25",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x3800
		x"70",x"F0",x"30",x"F0",x"F7",x"FF",x"F7",x"FF", -- 0x3808
		x"F7",x"FF",x"F7",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x3810
		x"F7",x"FF",x"F0",x"F0",x"F0",x"F0",x"80",x"00", -- 0x3818
		x"00",x"30",x"00",x"00",x"F0",x"C3",x"F0",x"F0", -- 0x3820
		x"F0",x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"FF", -- 0x3828
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF", -- 0x3830
		x"EF",x"FF",x"EF",x"FF",x"E7",x"FF",x"63",x"FF", -- 0x3838
		x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0", -- 0x3840
		x"70",x"F0",x"F7",x"FF",x"F7",x"FF",x"F7",x"FF", -- 0x3848
		x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3850
		x"F0",x"F1",x"F0",x"F0",x"00",x"00",x"00",x"00", -- 0x3858
		x"43",x"7F",x"73",x"FF",x"F3",x"FF",x"F7",x"FF", -- 0x3860
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3868
		x"FF",x"FF",x"DF",x"FF",x"DF",x"FF",x"DF",x"FF", -- 0x3870
		x"DF",x"FF",x"DF",x"FF",x"D7",x"FF",x"87",x"FF", -- 0x3878
		x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"F0",x"F1", -- 0x3880
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3888
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"F3", -- 0x3890
		x"F0",x"F1",x"00",x"10",x"00",x"10",x"00",x"10", -- 0x3898
		x"F7",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38A0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38A8
		x"BF",x"FF",x"BF",x"FF",x"BF",x"FF",x"BF",x"FF", -- 0x38B0
		x"BF",x"FF",x"BF",x"FF",x"1F",x"FF",x"FF",x"FF", -- 0x38B8
		x"F0",x"F0",x"F0",x"F1",x"F0",x"F3",x"FF",x"FF", -- 0x38C0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38D0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38D8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x38F8
		x"FF",x"E8",x"FF",x"E8",x"FF",x"E8",x"FF",x"E8", -- 0x3900
		x"FF",x"E8",x"FF",x"EC",x"FF",x"EC",x"FF",x"EC", -- 0x3908
		x"FF",x"EE",x"FF",x"EE",x"FF",x"FE",x"FF",x"FF", -- 0x3910
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3918
		x"00",x"30",x"00",x"31",x"00",x"31",x"00",x"31", -- 0x3920
		x"00",x"31",x"00",x"31",x"00",x"31",x"00",x"31", -- 0x3928
		x"00",x"31",x"00",x"31",x"00",x"31",x"00",x"31", -- 0x3930
		x"00",x"31",x"80",x"31",x"88",x"31",x"88",x"31", -- 0x3938
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3940
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3948
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3950
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3958
		x"CC",x"31",x"EC",x"31",x"FE",x"31",x"FF",x"F3", -- 0x3960
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3968
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3970
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3978
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3980
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3988
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3990
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3998
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A08
		x"FF",x"0F",x"8F",x"0F",x"8F",x"0F",x"0F",x"0F", -- 0x3A10
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3A18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A28
		x"7F",x"FF",x"1F",x"FF",x"1F",x"FF",x"0F",x"FF", -- 0x3A30
		x"0F",x"FF",x"0F",x"FF",x"0F",x"7F",x"0F",x"7F", -- 0x3A38
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3A40
		x"8F",x"0F",x"8F",x"0F",x"FF",x"0F",x"FF",x"FF", -- 0x3A48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A58
		x"0F",x"7F",x"0F",x"FF",x"0F",x"FF",x"0F",x"FF", -- 0x3A60
		x"0F",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3A98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"EF", -- 0x3AB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AD8
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3AF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B10
		x"FF",x"9F",x"FF",x"0F",x"EF",x"0F",x"EF",x"0F", -- 0x3B18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B30
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"7F",x"FF", -- 0x3B38
		x"EF",x"0F",x"FF",x"0F",x"FF",x"9F",x"FF",x"FF", -- 0x3B40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B58
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3B78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x3B80
		x"FF",x"0F",x"EF",x"0F",x"CF",x"0F",x"CF",x"0F", -- 0x3B88
		x"CF",x"0F",x"8F",x"0F",x"8F",x"0F",x"8F",x"0F", -- 0x3B90
		x"CF",x"0F",x"CF",x"0F",x"CF",x"0F",x"EF",x"0F", -- 0x3B98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x3BA0
		x"0F",x"FF",x"0F",x"7F",x"0F",x"3F",x"0F",x"3F", -- 0x3BA8
		x"0F",x"3F",x"0F",x"1F",x"0F",x"1F",x"0F",x"1F", -- 0x3BB0
		x"0F",x"3F",x"0F",x"3F",x"0F",x"7F",x"0F",x"7F", -- 0x3BB8
		x"FF",x"0F",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x3BC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BD8
		x"0F",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3BF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C38
		x"7F",x"FF",x"1F",x"FF",x"0F",x"FF",x"0F",x"FF", -- 0x3C40
		x"0F",x"FF",x"0F",x"FF",x"0F",x"FF",x"0F",x"FF", -- 0x3C48
		x"1F",x"FF",x"1F",x"FF",x"1F",x"FF",x"3F",x"FF", -- 0x3C50
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3C80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF", -- 0x3C88
		x"FF",x"CF",x"FF",x"8F",x"FF",x"8F",x"FF",x"8F", -- 0x3C90
		x"FF",x"CF",x"FF",x"CF",x"FF",x"EF",x"FF",x"FF", -- 0x3C98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF", -- 0x3CA8
		x"3F",x"FF",x"1F",x"FF",x"1F",x"FF",x"1F",x"FF", -- 0x3CB0
		x"1F",x"FF",x"1F",x"FF",x"3F",x"FF",x"8F",x"3F", -- 0x3CB8
		x"FF",x"FF",x"FF",x"EF",x"FF",x"EF",x"FF",x"EF", -- 0x3CC0
		x"FF",x"CF",x"FF",x"CF",x"FF",x"CF",x"FF",x"CF", -- 0x3CC8
		x"FF",x"EF",x"FF",x"EF",x"FF",x"EF",x"FF",x"FF", -- 0x3CD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3CD8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3CE0
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3CE8
		x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F", -- 0x3CF0
		x"8F",x"0F",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF", -- 0x3CF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D10
		x"FF",x"FF",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D30
		x"FF",x"FF",x"77",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF", -- 0x3D40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"FF", -- 0x3D60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3D98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F", -- 0x3DE0
		x"EF",x"1F",x"CF",x"0F",x"CF",x"0F",x"CF",x"0F", -- 0x3DE8
		x"EF",x"1F",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF", -- 0x3DF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E10
		x"FF",x"FF",x"FF",x"33",x"EE",x"DD",x"DD",x"EE", -- 0x3E18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E38
		x"DD",x"EE",x"DD",x"EE",x"EE",x"DD",x"FF",x"33", -- 0x3E40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EB0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3ED0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3ED8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3EF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"33",x"EE",x"DD", -- 0x3F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F20
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F38
		x"EE",x"DD",x"FF",x"33",x"FF",x"FF",x"FF",x"FF", -- 0x3F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F78
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3F88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"FF",x"CC", -- 0x3F90
		x"FF",x"DD",x"FF",x"CC",x"FF",x"EE",x"FF",x"FF", -- 0x3F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FA8
		x"FF",x"FF",x"FF",x"FF",x"33",x"FF",x"99",x"FF", -- 0x3FB0
		x"DD",x"FF",x"99",x"FF",x"33",x"FF",x"FF",x"FF", -- 0x3FB8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FC0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FD0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FD8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FE0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3FF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"  -- 0x3FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
