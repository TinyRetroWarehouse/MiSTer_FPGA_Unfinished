-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_A3 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_A3 is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"FB",x"FF",x"FF",x"FF",x"5F",x"0F",x"87",x"17", -- 0x0000
		x"CE",x"FD",x"5F",x"BF",x"FF",x"DD",x"CE",x"EE", -- 0x0008
		x"FF",x"FB",x"FF",x"FF",x"FF",x"BF",x"2F",x"87", -- 0x0010
		x"9B",x"9F",x"FF",x"FF",x"7F",x"DF",x"CF",x"67", -- 0x0018
		x"FE",x"FF",x"7F",x"9F",x"B7",x"99",x"DB",x"B1", -- 0x0020
		x"F8",x"B8",x"56",x"46",x"62",x"81",x"83",x"4F", -- 0x0028
		x"FF",x"FF",x"FF",x"F7",x"FF",x"FF",x"FD",x"FF", -- 0x0030
		x"FD",x"77",x"EC",x"C2",x"65",x"EF",x"A9",x"F3", -- 0x0038
		x"7F",x"BF",x"7A",x"F0",x"F9",x"AB",x"BB",x"97", -- 0x0040
		x"C7",x"E3",x"E3",x"49",x"F9",x"E2",x"77",x"BF", -- 0x0048
		x"FF",x"FF",x"FF",x"77",x"7B",x"FF",x"FF",x"FD", -- 0x0050
		x"FD",x"FF",x"FF",x"3F",x"1F",x"0F",x"09",x"CF", -- 0x0058
		x"FF",x"7F",x"7E",x"7F",x"FE",x"7C",x"5C",x"9E", -- 0x0060
		x"9E",x"BF",x"6F",x"37",x"12",x"1E",x"BE",x"EF", -- 0x0068
		x"FF",x"FF",x"F7",x"FF",x"FF",x"AD",x"1F",x"0F", -- 0x0070
		x"7D",x"FF",x"FF",x"FF",x"BF",x"1F",x"2F",x"7F", -- 0x0078
		x"FF",x"BF",x"FF",x"FF",x"4F",x"1F",x"1F",x"AF", -- 0x0080
		x"FF",x"BE",x"4C",x"5C",x"6E",x"97",x"8F",x"4F", -- 0x0088
		x"FF",x"DD",x"FD",x"FF",x"7F",x"7F",x"FB",x"F9", -- 0x0090
		x"BB",x"7F",x"1F",x"3F",x"1F",x"DF",x"FF",x"FF", -- 0x0098
		x"DF",x"B7",x"33",x"73",x"BF",x"5F",x"E7",x"E6", -- 0x00A0
		x"EA",x"A7",x"73",x"E2",x"E1",x"F5",x"DE",x"EE", -- 0x00A8
		x"FF",x"FF",x"FF",x"C7",x"CF",x"C7",x"63",x"F1", -- 0x00B0
		x"FB",x"FF",x"FF",x"FF",x"5F",x"FF",x"CF",x"E7", -- 0x00B8
		x"FF",x"FF",x"BF",x"BF",x"FB",x"F8",x"F0",x"F2", -- 0x00C0
		x"E9",x"FF",x"FF",x"F7",x"CF",x"E7",x"9E",x"EE", -- 0x00C8
		x"FF",x"FB",x"FB",x"FF",x"7F",x"FF",x"FF",x"7F", -- 0x00D0
		x"3F",x"F3",x"F7",x"E3",x"62",x"D5",x"DF",x"E7", -- 0x00D8
		x"FF",x"BE",x"FF",x"F7",x"FB",x"E7",x"E7",x"AF", -- 0x00E0
		x"DB",x"CB",x"E1",x"40",x"F0",x"E1",x"77",x"BF", -- 0x00E8
		x"FD",x"F7",x"E7",x"D9",x"DE",x"3F",x"8F",x"9F", -- 0x00F0
		x"CA",x"5D",x"17",x"0F",x"9B",x"86",x"89",x"CF", -- 0x00F8
		x"FF",x"9F",x"FD",x"FF",x"7F",x"FF",x"FF",x"DF", -- 0x0100
		x"FF",x"F8",x"E9",x"E8",x"DD",x"AF",x"3F",x"0F", -- 0x0108
		x"7F",x"BD",x"FB",x"E9",x"DE",x"87",x"8F",x"C5", -- 0x0110
		x"C0",x"E1",x"EF",x"DF",x"6F",x"76",x"09",x"CF", -- 0x0118
		x"FF",x"FF",x"FD",x"EB",x"80",x"C5",x"EF",x"EF", -- 0x0120
		x"D7",x"FF",x"FF",x"FF",x"FF",x"7E",x"74",x"F8", -- 0x0128
		x"FD",x"FB",x"FD",x"ED",x"CE",x"C7",x"C5",x"CA", -- 0x0130
		x"9A",x"B9",x"14",x"0A",x"2D",x"77",x"79",x"BB", -- 0x0138
		x"FB",x"DD",x"FF",x"FF",x"EF",x"FE",x"9E",x"8F", -- 0x0140
		x"1F",x"0F",x"03",x"03",x"9F",x"FF",x"EF",x"FC", -- 0x0148
		x"FF",x"FB",x"F9",x"DD",x"2F",x"1F",x"0F",x"7F", -- 0x0150
		x"FE",x"DD",x"F0",x"EA",x"DD",x"9F",x"09",x"1B", -- 0x0158
		x"FF",x"DE",x"BE",x"FE",x"FF",x"FF",x"F7",x"E7", -- 0x0160
		x"EE",x"C7",x"CB",x"C2",x"A1",x"E2",x"7E",x"2E", -- 0x0168
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"15",x"8B", -- 0x0170
		x"C7",x"E7",x"B7",x"D3",x"62",x"D5",x"DF",x"E7", -- 0x0178
		x"9F",x"C3",x"65",x"CF",x"C7",x"8B",x"47",x"2F", -- 0x0180
		x"3F",x"FF",x"FB",x"B3",x"F1",x"F8",x"E9",x"FF", -- 0x0188
		x"CE",x"B3",x"13",x"9F",x"BF",x"FF",x"FF",x"DF", -- 0x0190
		x"9F",x"8F",x"DF",x"FF",x"FF",x"FD",x"FF",x"FF", -- 0x0198
		x"1F",x"8F",x"6C",x"F1",x"FC",x"AD",x"B1",x"98", -- 0x01A0
		x"D8",x"FE",x"FE",x"57",x"EF",x"7F",x"3F",x"7F", -- 0x01A8
		x"EF",x"AB",x"E3",x"71",x"70",x"39",x"89",x"DC", -- 0x01B0
		x"C9",x"1D",x"1F",x"0B",x"07",x"0F",x"FF",x"FF", -- 0x01B8
		x"2E",x"47",x"17",x"1C",x"DD",x"79",x"79",x"38", -- 0x01C0
		x"98",x"FC",x"6F",x"3E",x"7C",x"7C",x"3C",x"7F", -- 0x01C8
		x"19",x"3F",x"3F",x"97",x"8F",x"9F",x"7D",x"FF", -- 0x01D0
		x"7F",x"7F",x"FF",x"DF",x"1F",x"4F",x"6F",x"7F", -- 0x01D8
		x"EF",x"47",x"02",x"01",x"C3",x"72",x"7A",x"BF", -- 0x01E0
		x"9F",x"DF",x"67",x"3F",x"7E",x"2C",x"9C",x"BE", -- 0x01E8
		x"FF",x"FF",x"FF",x"EF",x"5F",x"1F",x"6F",x"3F", -- 0x01F0
		x"FF",x"FF",x"7F",x"FF",x"BD",x"1D",x"4F",x"7F", -- 0x01F8
		x"EE",x"47",x"07",x"43",x"E3",x"77",x"2F",x"3E", -- 0x0200
		x"3E",x"6F",x"E7",x"C3",x"C7",x"EE",x"BC",x"FC", -- 0x0208
		x"FF",x"FB",x"FF",x"FF",x"BF",x"5F",x"0D",x"1F", -- 0x0210
		x"1F",x"3F",x"FF",x"FD",x"FD",x"7F",x"3F",x"7F", -- 0x0218
		x"1F",x"97",x"72",x"F2",x"F1",x"BB",x"BF",x"9D", -- 0x0220
		x"D3",x"C3",x"E7",x"4D",x"E5",x"E0",x"75",x"BE", -- 0x0228
		x"C4",x"A1",x"13",x"1F",x"3F",x"1F",x"8F",x"CF", -- 0x0230
		x"EF",x"7F",x"FB",x"FF",x"3F",x"3F",x"7D",x"EF", -- 0x0238
		x"3F",x"1F",x"8D",x"83",x"C6",x"C0",x"E2",x"BF", -- 0x0240
		x"FF",x"DF",x"FF",x"EF",x"C2",x"C9",x"FF",x"FF", -- 0x0248
		x"F7",x"AB",x"D3",x"E1",x"52",x"05",x"0F",x"06", -- 0x0250
		x"C2",x"C1",x"E7",x"FF",x"EF",x"FF",x"FB",x"FF", -- 0x0258
		x"EE",x"47",x"05",x"00",x"C0",x"72",x"7D",x"3F", -- 0x0260
		x"09",x"38",x"F0",x"B9",x"FF",x"EE",x"E4",x"FC", -- 0x0268
		x"19",x"BE",x"FF",x"DF",x"17",x"06",x"C4",x"D0", -- 0x0270
		x"5C",x"06",x"0E",x"83",x"C3",x"65",x"E0",x"70", -- 0x0278
		x"4F",x"26",x"A7",x"C0",x"F0",x"DE",x"AE",x"18", -- 0x0280
		x"1A",x"8E",x"CC",x"5E",x"8F",x"07",x"AF",x"FF", -- 0x0288
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"D5",x"6B", -- 0x0290
		x"FF",x"57",x"37",x"03",x"82",x"D1",x"F8",x"FC", -- 0x0298
		x"FF",x"BE",x"FF",x"F7",x"FF",x"FF",x"F9",x"D0", -- 0x02A0
		x"E3",x"F3",x"F1",x"B8",x"BC",x"FC",x"F9",x"FF", -- 0x02A8
		x"17",x"4B",x"53",x"21",x"22",x"C1",x"F7",x"E1", -- 0x02B0
		x"E0",x"79",x"F9",x"F1",x"F8",x"F8",x"FC",x"FC", -- 0x02B8
		x"FE",x"BE",x"9F",x"BF",x"FF",x"F7",x"E7",x"E3", -- 0x02C0
		x"E7",x"FE",x"FD",x"A9",x"F8",x"D0",x"F9",x"FF", -- 0x02C8
		x"49",x"33",x"15",x"C1",x"C2",x"E3",x"F1",x"FC", -- 0x02D0
		x"FD",x"BF",x"DF",x"8F",x"87",x"BF",x"FD",x"FF", -- 0x02D8
		x"5F",x"3E",x"37",x"A4",x"CC",x"8E",x"C7",x"E7", -- 0x02E0
		x"EF",x"C5",x"C3",x"E3",x"C1",x"F0",x"F8",x"FE", -- 0x02E8
		x"5F",x"67",x"2B",x"3F",x"5F",x"15",x"01",x"9B", -- 0x02F0
		x"FF",x"D7",x"C7",x"E3",x"BA",x"5D",x"5F",x"27", -- 0x02F8
		x"FE",x"FC",x"99",x"D8",x"F3",x"F0",x"F8",x"F8", -- 0x0300
		x"BF",x"BE",x"FE",x"FE",x"EC",x"FC",x"BC",x"FA", -- 0x0308
		x"5F",x"E7",x"EB",x"DF",x"CF",x"C5",x"45",x"CB", -- 0x0310
		x"1F",x"77",x"77",x"93",x"62",x"75",x"5F",x"27", -- 0x0318
		x"DF",x"BF",x"35",x"74",x"B9",x"56",x"EE",x"F6", -- 0x0320
		x"C4",x"84",x"6A",x"F2",x"F1",x"E1",x"DC",x"ED", -- 0x0328
		x"FF",x"FF",x"77",x"FF",x"7F",x"FF",x"79",x"FD", -- 0x0330
		x"7F",x"3F",x"FF",x"EF",x"6F",x"7B",x"FF",x"FF", -- 0x0338
		x"EE",x"4F",x"13",x"10",x"C1",x"79",x"3D",x"1E", -- 0x0340
		x"13",x"B0",x"F9",x"FF",x"FF",x"BE",x"9F",x"FF", -- 0x0348
		x"19",x"3E",x"3F",x"DF",x"D7",x"EA",x"C0",x"C0", -- 0x0350
		x"EE",x"FF",x"FF",x"FF",x"7B",x"FB",x"FF",x"FF", -- 0x0358
		x"FF",x"DF",x"BD",x"FD",x"FF",x"FF",x"EE",x"C6", -- 0x0360
		x"CE",x"E6",x"E6",x"F3",x"7F",x"7B",x"BA",x"ED", -- 0x0368
		x"FF",x"EF",x"FF",x"FB",x"FF",x"3F",x"FF",x"7F", -- 0x0370
		x"5B",x"33",x"02",x"51",x"13",x"B9",x"74",x"7E", -- 0x0378
		x"FF",x"BD",x"E9",x"DF",x"8D",x"1F",x"0B",x"07", -- 0x0380
		x"8B",x"81",x"C6",x"EF",x"CB",x"C7",x"93",x"CF", -- 0x0388
		x"FF",x"FF",x"FF",x"DB",x"D9",x"FF",x"FF",x"FF", -- 0x0390
		x"EF",x"7F",x"FF",x"FF",x"D7",x"8F",x"07",x"8F", -- 0x0398
		x"BF",x"DD",x"FF",x"FB",x"F1",x"70",x"F1",x"F9", -- 0x03A0
		x"EF",x"C6",x"CF",x"FF",x"FB",x"BC",x"BF",x"FF", -- 0x03A8
		x"FF",x"F7",x"FB",x"DF",x"8B",x"07",x"0F",x"05", -- 0x03B0
		x"03",x"83",x"DF",x"FF",x"EF",x"C3",x"C7",x"FF", -- 0x03B8
		x"EE",x"47",x"07",x"01",x"C3",x"70",x"79",x"3B", -- 0x03C0
		x"01",x"00",x"00",x"00",x"62",x"A0",x"B5",x"D7", -- 0x03C8
		x"19",x"3E",x"3F",x"DF",x"57",x"E6",x"E4",x"F0", -- 0x03D0
		x"5C",x"06",x"0E",x"03",x"03",x"05",x"00",x"20", -- 0x03D8
		x"3F",x"1F",x"0C",x"03",x"06",x"00",x"00",x"04", -- 0x03E0
		x"A4",x"AA",x"AA",x"9B",x"91",x"B9",x"AA",x"4A", -- 0x03E8
		x"F7",x"AB",x"13",x"21",x"12",x"05",x"0F",x"06", -- 0x03F0
		x"02",x"00",x"01",x"0B",x"0D",x"6C",x"64",x"42", -- 0x03F8
		x"EE",x"47",x"07",x"01",x"C3",x"70",x"39",x"1F", -- 0x0400
		x"03",x"00",x"80",x"80",x"A3",x"63",x"6B",x"49", -- 0x0408
		x"19",x"3E",x"3F",x"DF",x"57",x"EA",x"C0",x"80", -- 0x0410
		x"80",x"80",x"A2",x"FE",x"5A",x"49",x"65",x"35", -- 0x0418
		x"9F",x"C3",x"6D",x"9F",x"97",x"8E",x"40",x"20", -- 0x0420
		x"0D",x"0D",x"2D",x"A4",x"2A",x"AA",x"AA",x"95", -- 0x0428
		x"CE",x"B2",x"31",x"81",x"01",x"95",x"96",x"3A", -- 0x0430
		x"2A",x"3A",x"51",x"55",x"C5",x"A5",x"AA",x"22", -- 0x0438
		x"DF",x"BE",x"37",x"74",x"B8",x"56",x"EF",x"F6", -- 0x0440
		x"EE",x"A7",x"43",x"82",x"C1",x"E5",x"DE",x"EE", -- 0x0448
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"D5",x"EB", -- 0x0450
		x"FF",x"77",x"77",x"D3",x"62",x"D5",x"DF",x"E7", -- 0x0458
		x"9D",x"DB",x"6D",x"9E",x"B5",x"9F",x"D9",x"A6", -- 0x0460
		x"77",x"BA",x"50",x"54",x"66",x"99",x"87",x"4F", -- 0x0468
		x"C9",x"B3",x"2D",x"CD",x"8E",x"C7",x"65",x"42", -- 0x0470
		x"2A",x"71",x"D4",x"4A",x"6D",x"37",x"19",x"BB", -- 0x0478
		x"3F",x"9F",x"6C",x"F3",x"FA",x"AD",x"B3",x"97", -- 0x0480
		x"DF",x"C5",x"E1",x"4C",x"F0",x"E2",x"77",x"BF", -- 0x0488
		x"F7",x"AB",x"D3",x"61",x"52",x"05",x"8F",x"DF", -- 0x0490
		x"EA",x"5D",x"1F",x"2F",x"1B",x"06",x"09",x"CF", -- 0x0498
		x"EE",x"47",x"07",x"01",x"C3",x"70",x"79",x"BF", -- 0x04A0
		x"93",x"F8",x"69",x"36",x"72",x"3E",x"BF",x"EF", -- 0x04A8
		x"19",x"3E",x"3F",x"DF",x"57",x"E6",x"E4",x"F0", -- 0x04B0
		x"7C",x"D6",x"E6",x"F3",x"E3",x"79",x"34",x"FE", -- 0x04B8
		x"00",x"02",x"20",x"00",x"00",x"02",x"00",x"00", -- 0x04C0
		x"00",x"00",x"00",x"20",x"00",x"00",x"01",x"00", -- 0x04C8
		x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00", -- 0x04D0
		x"00",x"00",x"00",x"00",x"82",x"40",x"00",x"00", -- 0x04D8
		x"00",x"08",x"48",x"00",x"09",x"20",x"00",x"00", -- 0x04E0
		x"00",x"00",x"02",x"18",x"00",x"00",x"00",x"00", -- 0x04E8
		x"00",x"00",x"04",x"08",x"08",x"00",x"20",x"50", -- 0x04F0
		x"00",x"04",x"02",x"16",x"10",x"30",x"08",x"00", -- 0x04F8
		x"DF",x"ED",x"FB",x"BB",x"DE",x"FB",x"B1",x"BE", -- 0x0500
		x"FD",x"D8",x"FE",x"EF",x"EE",x"BD",x"9E",x"FF", -- 0x0508
		x"00",x"30",x"20",x"60",x"40",x"40",x"2C",x"46", -- 0x0510
		x"C2",x"1D",x"97",x"8B",x"99",x"F3",x"AE",x"FF", -- 0x0518
		x"80",x"80",x"20",x"C0",x"88",x"5C",x"88",x"91", -- 0x0520
		x"D9",x"AE",x"FF",x"AF",x"F6",x"E7",x"71",x"FF", -- 0x0528
		x"00",x"00",x"00",x"10",x"20",x"70",x"20",x"E8", -- 0x0530
		x"46",x"C3",x"87",x"85",x"ED",x"AD",x"97",x"FF", -- 0x0538
		x"80",x"80",x"C0",x"D8",x"F0",x"A1",x"66",x"CE", -- 0x0540
		x"FD",x"94",x"C8",x"DB",x"E9",x"F1",x"EE",x"FF", -- 0x0548
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"50", -- 0x0550
		x"20",x"C0",x"A0",x"60",x"24",x"18",x"BC",x"EF", -- 0x0558
		x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"08", -- 0x0560
		x"A8",x"DC",x"86",x"86",x"DD",x"FA",x"A7",x"FF", -- 0x0568
		x"00",x"00",x"40",x"20",x"30",x"18",x"10",x"00", -- 0x0570
		x"00",x"00",x"00",x"C0",x"60",x"E0",x"98",x"FE", -- 0x0578
		x"80",x"C0",x"C0",x"A0",x"E0",x"B8",x"A0",x"D0", -- 0x0580
		x"D0",x"F0",x"49",x"9A",x"86",x"DE",x"B9",x"FD", -- 0x0588
		x"00",x"20",x"50",x"38",x"20",x"00",x"00",x"00", -- 0x0590
		x"00",x"40",x"10",x"20",x"00",x"00",x"00",x"00", -- 0x0598
		x"00",x"00",x"04",x"03",x"0B",x"02",x"04",x"80", -- 0x05A0
		x"80",x"E2",x"C2",x"84",x"38",x"48",x"8D",x"FE", -- 0x05A8
		x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"20", -- 0x05B0
		x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05B8
		x"BE",x"F8",x"D9",x"B7",x"7D",x"B0",x"E3",x"DF", -- 0x05C0
		x"FD",x"F4",x"CE",x"D9",x"6B",x"ED",x"DE",x"7F", -- 0x05C8
		x"00",x"00",x"80",x"00",x"A0",x"C0",x"A0",x"D0", -- 0x05D0
		x"80",x"04",x"32",x"36",x"9C",x"F4",x"AC",x"9F", -- 0x05D8
		x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x05E0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05E8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x05F8
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF", -- 0x0600
		x"FF",x"FF",x"FF",x"DF",x"FB",x"FF",x"FF",x"FF", -- 0x0608
		x"FF",x"EF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FB", -- 0x0610
		x"F7",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x0618
		x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"DF",x"FF", -- 0x0620
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0628
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0630
		x"FF",x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x0638
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0640
		x"FF",x"FE",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF", -- 0x0648
		x"FF",x"FF",x"FF",x"FF",x"BF",x"FF",x"FF",x"FF", -- 0x0650
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0658
		x"FF",x"F7",x"DF",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x0660
		x"EF",x"63",x"97",x"87",x"83",x"09",x"09",x"BF", -- 0x0668
		x"FF",x"F7",x"FF",x"3F",x"FF",x"FF",x"FF",x"FF", -- 0x0670
		x"FB",x"FB",x"FF",x"BF",x"FF",x"FD",x"FF",x"FF", -- 0x0678
		x"FF",x"EF",x"EF",x"FF",x"FF",x"FF",x"BF",x"FF", -- 0x0680
		x"FD",x"FF",x"FE",x"AC",x"B0",x"F8",x"FC",x"FC", -- 0x0688
		x"FF",x"FF",x"E7",x"FF",x"BF",x"FF",x"FF",x"FF", -- 0x0690
		x"BF",x"D7",x"EF",x"27",x"0F",x"25",x"73",x"3F", -- 0x0698
		x"00",x"02",x"03",x"03",x"07",x"01",x"02",x"01", -- 0x06A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06A8
		x"00",x"00",x"00",x"80",x"80",x"C0",x"00",x"80", -- 0x06B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C8
		x"00",x"18",x"1C",x"0C",x"1C",x"14",x"08",x"00", -- 0x06D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06D8
		x"00",x"40",x"00",x"02",x"00",x"08",x"0B",x"00", -- 0x06E0
		x"30",x"00",x"04",x"04",x"40",x"00",x"00",x"00", -- 0x06E8
		x"00",x"20",x"30",x"20",x"00",x"80",x"80",x"04", -- 0x06F0
		x"00",x"00",x"00",x"08",x"12",x"04",x"10",x"00", -- 0x06F8
		x"00",x"04",x"02",x"04",x"00",x"00",x"04",x"30", -- 0x0700
		x"B1",x"B3",x"77",x"AF",x"F2",x"C9",x"30",x"F1", -- 0x0708
		x"00",x"00",x"08",x"00",x"00",x"00",x"10",x"CA", -- 0x0710
		x"67",x"41",x"13",x"98",x"8C",x"8F",x"F7",x"FF", -- 0x0718
		x"00",x"01",x"02",x"00",x"10",x"00",x"01",x"03", -- 0x0720
		x"01",x"01",x"00",x"08",x"1C",x"0E",x"02",x"10", -- 0x0728
		x"F7",x"B3",x"F9",x"8F",x"2D",x"31",x"31",x"B0", -- 0x0730
		x"84",x"FB",x"BF",x"3D",x"39",x"23",x"72",x"DF", -- 0x0738
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0740
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0748
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0750
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0760
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0768
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0770
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0778
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0798
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F8
		x"90",x"80",x"74",x"68",x"24",x"A0",x"D0",x"54", -- 0x0800
		x"4A",x"EA",x"A4",x"36",x"74",x"59",x"1E",x"A7", -- 0x0808
		x"F7",x"FB",x"7F",x"7F",x"3F",x"3F",x"3F",x"3D", -- 0x0810
		x"1F",x"1F",x"0F",x"87",x"07",x"03",x"43",x"21", -- 0x0818
		x"FF",x"7F",x"3F",x"3F",x"1F",x"0F",x"47",x"07", -- 0x0820
		x"83",x"43",x"83",x"51",x"A0",x"50",x"D0",x"A4", -- 0x0828
		x"FF",x"F7",x"FB",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x0830
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x0838
		x"40",x"21",x"89",x"01",x"50",x"90",x"08",x"A0", -- 0x0840
		x"A0",x"44",x"50",x"48",x"E0",x"A0",x"28",x"10", -- 0x0848
		x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x0850
		x"7F",x"FF",x"FD",x"7D",x"7F",x"FF",x"FF",x"FF", -- 0x0858
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0860
		x"3F",x"0D",x"00",x"00",x"A0",x"14",x"01",x"AA", -- 0x0868
		x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"7F",x"BF", -- 0x0870
		x"FF",x"FF",x"EF",x"FF",x"7F",x"1F",x"03",x"41", -- 0x0878
		x"FF",x"FF",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0880
		x"3F",x"0F",x"83",x"81",x"31",x"80",x"48",x"B0", -- 0x0888
		x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD", -- 0x0890
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0898
		x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"9C", -- 0x08A0
		x"00",x"00",x"12",x"26",x"98",x"65",x"AA",x"59", -- 0x08A8
		x"FF",x"FF",x"FF",x"DF",x"7F",x"FF",x"7F",x"FF", -- 0x08B0
		x"3C",x"00",x"00",x"82",x"20",x"48",x"05",x"AA", -- 0x08B8
		x"FF",x"3F",x"13",x"01",x"01",x"40",x"02",x"D0", -- 0x08C0
		x"24",x"B5",x"A8",x"4A",x"52",x"37",x"99",x"4A", -- 0x08C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"07",x"03", -- 0x08D0
		x"00",x"40",x"20",x"8A",x"D0",x"2A",x"01",x"AD", -- 0x08D8
		x"90",x"80",x"A8",x"72",x"40",x"D4",x"69",x"DC", -- 0x08E0
		x"CA",x"AB",x"B5",x"D5",x"55",x"7A",x"2A",x"A5", -- 0x08E8
		x"FF",x"7F",x"6F",x"1F",x"1F",x"0F",x"03",x"41", -- 0x08F0
		x"A0",x"80",x"50",x"A4",x"95",x"58",x"AA",x"2B", -- 0x08F8
		x"FF",x"7F",x"2F",x"07",x"07",x"43",x"02",x"A1", -- 0x0900
		x"41",x"10",x"A0",x"10",x"A8",x"6D",x"49",x"B2", -- 0x0908
		x"FF",x"FF",x"FF",x"FB",x"F9",x"FF",x"FF",x"FF", -- 0x0910
		x"DF",x"9F",x"2F",x"1F",x"0F",x"03",x"03",x"41", -- 0x0918
		x"29",x"69",x"B2",x"14",x"60",x"8A",x"39",x"A9", -- 0x0920
		x"C5",x"1F",x"51",x"03",x"2A",x"B5",x"58",x"39", -- 0x0928
		x"80",x"50",x"00",x"AA",x"A4",x"B5",x"70",x"52", -- 0x0930
		x"49",x"29",x"A0",x"32",x"50",x"1D",x"54",x"66", -- 0x0938
		x"66",x"2A",x"B8",x"0A",x"4C",x"05",x"95",x"B2", -- 0x0940
		x"4A",x"AE",x"AF",x"A5",x"95",x"D1",x"CA",x"29", -- 0x0948
		x"FC",x"3A",x"AD",x"55",x"C1",x"AA",x"F8",x"A3", -- 0x0950
		x"95",x"9F",x"51",x"06",x"A8",x"CD",x"96",x"94", -- 0x0958
		x"29",x"69",x"B2",x"14",x"60",x"8A",x"39",x"A9", -- 0x0960
		x"C5",x"1F",x"51",x"03",x"2A",x"B5",x"58",x"39", -- 0x0968
		x"94",x"52",x"02",x"A8",x"A5",x"B5",x"70",x"52", -- 0x0970
		x"49",x"29",x"A0",x"32",x"50",x"1D",x"54",x"66", -- 0x0978
		x"FF",x"7F",x"7F",x"3F",x"1F",x"3F",x"3F",x"3F", -- 0x0980
		x"1F",x"1F",x"9D",x"0F",x"0F",x"0F",x"8F",x"8F", -- 0x0988
		x"FF",x"F7",x"FB",x"F7",x"FF",x"FF",x"FF",x"FF", -- 0x0990
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x0998
		x"0F",x"0F",x"8F",x"05",x"43",x"83",x"03",x"A3", -- 0x09A0
		x"A1",x"43",x"43",x"41",x"E0",x"A0",x"28",x"10", -- 0x09A8
		x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x09B0
		x"FF",x"FF",x"FD",x"7D",x"7F",x"FF",x"FF",x"FF", -- 0x09B8
		x"90",x"80",x"74",x"68",x"24",x"A0",x"D0",x"54", -- 0x09C0
		x"4A",x"EA",x"A4",x"36",x"74",x"59",x"1E",x"A7", -- 0x09C8
		x"F7",x"FB",x"7F",x"7F",x"7F",x"3F",x"3F",x"3D", -- 0x09D0
		x"3F",x"3F",x"1F",x"9F",x"0F",x"0F",x"4F",x"0F", -- 0x09D8
		x"91",x"80",x"74",x"6A",x"25",x"A1",x"D1",x"54", -- 0x09E0
		x"4A",x"EA",x"A4",x"36",x"74",x"D9",x"5E",x"27", -- 0x09E8
		x"07",x"8B",x"87",x"07",x"47",x"47",x"25",x"A3", -- 0x09F0
		x"83",x"C3",x"13",x"83",x"61",x"21",x"51",x"21", -- 0x09F8
		x"0F",x"8F",x"87",x"03",x"23",x"41",x"00",x"A0", -- 0x0A00
		x"40",x"14",x"A4",x"11",x"A8",x"6D",x"49",x"B2", -- 0x0A08
		x"FF",x"FF",x"FF",x"FB",x"F9",x"FF",x"FF",x"FF", -- 0x0A10
		x"DF",x"1F",x"2F",x"1F",x"0F",x"03",x"03",x"51", -- 0x0A18
		x"40",x"22",x"88",x"02",x"52",x"90",x"08",x"A2", -- 0x0A20
		x"A0",x"44",x"51",x"49",x"E0",x"A0",x"28",x"10", -- 0x0A28
		x"8F",x"0F",x"8B",x"1F",x"1F",x"1F",x"9F",x"8F", -- 0x0A30
		x"07",x"07",x"0D",x"1D",x"1F",x"1F",x"8F",x"0F", -- 0x0A38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0A58
		x"C7",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC", -- 0x0A60
		x"FC",x"FC",x"FC",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x0A68
		x"07",x"07",x"0F",x"08",x"00",x"00",x"00",x"10", -- 0x0A70
		x"11",x"13",x"03",x"03",x"07",x"3F",x"3F",x"3F", -- 0x0A78
		x"D9",x"57",x"B7",x"F1",x"4D",x"FE",x"9D",x"DC", -- 0x0A80
		x"3A",x"C8",x"B2",x"92",x"0E",x"AB",x"21",x"A3", -- 0x0A88
		x"94",x"EA",x"72",x"CC",x"B4",x"D6",x"FF",x"FF", -- 0x0A90
		x"FF",x"FF",x"07",x"07",x"D7",x"90",x"28",x"54", -- 0x0A98
		x"55",x"73",x"FA",x"C8",x"E9",x"CF",x"EF",x"CA", -- 0x0AA0
		x"E9",x"FC",x"FE",x"FD",x"FE",x"FE",x"07",x"54", -- 0x0AA8
		x"A8",x"67",x"87",x"D7",x"F7",x"57",x"77",x"A7", -- 0x0AB0
		x"A7",x"57",x"C7",x"77",x"A7",x"E7",x"F0",x"B4", -- 0x0AB8
		x"55",x"73",x"FA",x"CF",x"AF",x"CF",x"66",x"46", -- 0x0AC0
		x"A7",x"76",x"A6",x"A1",x"D6",x"6A",x"FF",x"54", -- 0x0AC8
		x"A8",x"67",x"87",x"FF",x"FF",x"FF",x"07",x"A7", -- 0x0AD0
		x"A7",x"57",x"C7",x"77",x"A7",x"E7",x"F0",x"B4", -- 0x0AD8
		x"DB",x"BD",x"FF",x"A6",x"45",x"7F",x"75",x"6F", -- 0x0AE0
		x"45",x"43",x"47",x"00",x"A5",x"DB",x"57",x"54", -- 0x0AE8
		x"30",x"9F",x"9F",x"DF",x"1F",x"FF",x"FF",x"FF", -- 0x0AF0
		x"FF",x"FF",x"FF",x"1F",x"1F",x"00",x"90",x"DC", -- 0x0AF8
		x"BA",x"97",x"B7",x"F1",x"4D",x"EE",x"8D",x"4D", -- 0x0B00
		x"AE",x"CD",x"BF",x"3F",x"3F",x"80",x"21",x"A3", -- 0x0B08
		x"A4",x"E9",x"71",x"C9",x"B5",x"D1",x"6F",x"CF", -- 0x0B10
		x"8F",x"2F",x"FF",x"FF",x"FF",x"00",x"28",x"54", -- 0x0B18
		x"FF",x"C7",x"97",x"93",x"93",x"83",x"8B",x"F8", -- 0x0B20
		x"FF",x"FF",x"BF",x"BF",x"BF",x"83",x"FF",x"FF", -- 0x0B28
		x"FF",x"E1",x"DF",x"C1",x"C1",x"C1",x"DF",x"C1", -- 0x0B30
		x"C1",x"C1",x"DF",x"C1",x"C1",x"C3",x"FF",x"FF", -- 0x0B38
		x"FF",x"FF",x"BB",x"BB",x"9B",x"F8",x"C0",x"BF", -- 0x0B40
		x"80",x"80",x"81",x"E4",x"C4",x"C4",x"C4",x"C0", -- 0x0B48
		x"FF",x"E1",x"DF",x"C1",x"C1",x"C3",x"FF",x"FF", -- 0x0B50
		x"7F",x"7F",x"0F",x"5F",x"4F",x"4F",x"43",x"3F", -- 0x0B58
		x"FF",x"E1",x"DF",x"C1",x"C1",x"C1",x"DF",x"C1", -- 0x0B60
		x"C1",x"C3",x"FF",x"F0",x"EF",x"E0",x"E0",x"E0", -- 0x0B68
		x"FF",x"FF",x"7F",x"7F",x"7F",x"77",x"77",x"77", -- 0x0B70
		x"17",x"F3",x"E3",x"5F",x"C3",x"43",x"47",x"FF", -- 0x0B78
		x"FF",x"C3",x"BF",x"83",x"87",x"FF",x"FF",x"F7", -- 0x0B80
		x"E7",x"E3",x"E1",x"F3",x"FF",x"83",x"87",x"FF", -- 0x0B88
		x"FF",x"FF",x"FF",x"DF",x"9F",x"8F",x"87",x"CF", -- 0x0B90
		x"FF",x"FF",x"FF",x"BF",x"3F",x"1F",x"0F",x"9F", -- 0x0B98
		x"00",x"4A",x"AE",x"57",x"D5",x"2B",x"53",x"D5", -- 0x0BA0
		x"2B",x"55",x"B7",x"AC",x"D2",x"6D",x"25",x"D4", -- 0x0BA8
		x"00",x"14",x"B7",x"AB",x"7C",x"77",x"BB",x"AA", -- 0x0BB0
		x"65",x"7D",x"DE",x"AA",x"DB",x"56",x"55",x"AA", -- 0x0BB8
		x"EB",x"AE",x"77",x"55",x"5E",x"FB",x"AA",x"AE", -- 0x0BC0
		x"A5",x"EE",x"7A",x"5A",x"D7",x"BD",x"ED",x"ED", -- 0x0BC8
		x"34",x"AC",x"AA",x"88",x"5C",x"F4",x"BE",x"D4", -- 0x0BD0
		x"AC",x"FC",x"AC",x"F8",x"56",x"74",x"F4",x"6A", -- 0x0BD8
		x"00",x"22",x"67",x"55",x"5E",x"FB",x"AA",x"AE", -- 0x0BE0
		x"A5",x"EE",x"7A",x"5A",x"D7",x"BD",x"ED",x"ED", -- 0x0BE8
		x"00",x"00",x"A8",x"8A",x"5C",x"F4",x"BE",x"D6", -- 0x0BF0
		x"AC",x"FC",x"AC",x"F8",x"54",x"74",x"F6",x"68", -- 0x0BF8
		x"5F",x"BE",x"F7",x"54",x"68",x"1E",x"2F",x"96", -- 0x0C00
		x"8E",x"C7",x"43",x"61",x"38",x"39",x"12",x"11", -- 0x0C08
		x"5F",x"67",x"2B",x"3F",x"5F",x"3D",x"D5",x"EB", -- 0x0C10
		x"FF",x"77",x"77",x"D3",x"62",x"F5",x"FF",x"27", -- 0x0C18
		x"0C",x"0C",x"66",x"73",x"61",x"00",x"03",x"06", -- 0x0C20
		x"0C",x"3E",x"FC",x"D9",x"87",x"09",x"79",x"F0", -- 0x0C28
		x"77",x"3B",x"53",x"09",x"82",x"C1",x"67",x"65", -- 0x0C30
		x"62",x"CF",x"D4",x"8A",x"2D",x"3F",x"99",x"9B", -- 0x0C38
		x"31",x"00",x"00",x"01",x"00",x"08",x"08",x"90", -- 0x0C40
		x"E0",x"41",x"07",x"1C",x"30",x"C0",x"20",x"98", -- 0x0C48
		x"97",x"DB",x"B3",x"81",x"C2",x"C1",x"67",x"61", -- 0x0C50
		x"C2",x"61",x"31",x"31",x"18",x"19",x"18",x"0C", -- 0x0C58
		x"3F",x"1F",x"8D",x"40",x"22",x"1F",x"09",x"80", -- 0x0C60
		x"E0",x"C2",x"C2",x"64",x"20",x"20",x"01",x"43", -- 0x0C68
		x"F7",x"AB",x"D3",x"E1",x"52",x"45",x"07",x"82", -- 0x0C70
		x"59",x"2D",x"06",x"00",x"00",x"00",x"80",x"00", -- 0x0C78
		x"6F",x"CF",x"9E",x"9C",x"00",x"0C",x"0F",x"7E", -- 0x0C80
		x"78",x"F0",x"60",x"41",x"43",x"9F",x"3E",x"78", -- 0x0C88
		x"86",x"0C",x"0C",x"18",x"3C",x"78",x"B0",x"20", -- 0x0C90
		x"20",x"E1",x"C3",x"C7",x"C7",x"8E",x"1E",x"08", -- 0x0C98
		x"80",x"03",x"36",x"CC",x"31",x"0E",x"03",x"00", -- 0x0CA0
		x"00",x"02",x"01",x"00",x"C0",x"E3",x"FF",x"FF", -- 0x0CA8
		x"40",x"00",x"63",x"FE",x"9E",x"8C",x"40",x"30", -- 0x0CB0
		x"1F",x"03",x"C0",x"20",x"1B",x"86",x"E0",x"FF", -- 0x0CB8
		x"FE",x"BC",x"FE",x"F4",x"FC",x"FE",x"FF",x"DF", -- 0x0CC0
		x"EF",x"FF",x"FF",x"BF",x"BF",x"F3",x"C1",x"21", -- 0x0CC8
		x"17",x"4B",x"13",x"01",x"02",x"81",x"87",x"C1", -- 0x0CD0
		x"82",x"C1",x"D1",x"E1",x"E0",x"70",x"18",x"04", -- 0x0CD8
		x"F1",x"78",x"38",x"39",x"3C",x"1C",x"9C",x"CE", -- 0x0CE0
		x"CE",x"C7",x"E7",x"67",x"13",x"13",x"C3",x"E1", -- 0x0CE8
		x"00",x"80",x"C8",x"CC",x"CC",x"9C",x"9C",x"49", -- 0x0CF0
		x"48",x"4C",x"64",x"72",x"B3",x"B3",x"B9",x"D9", -- 0x0CF8
		x"71",x"79",x"3C",x"3C",x"19",x"19",x"09",x"8C", -- 0x0D00
		x"86",x"C7",x"E3",x"E3",x"F1",x"71",x"38",x"1C", -- 0x0D08
		x"83",x"C2",x"84",x"45",x"8D",x"8B",x"C7",x"E7", -- 0x0D10
		x"E6",x"66",x"63",x"33",x"B2",x"B8",x"D9",x"D9", -- 0x0D18
		x"0C",x"06",x"07",x"02",x"00",x"40",x"E0",x"F0", -- 0x0D20
		x"40",x"B3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D28
		x"16",x"0D",x"4A",x"00",x"02",x"00",x"00",x"02", -- 0x0D30
		x"C0",x"3A",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D38
		x"00",x"01",x"02",x"00",x"10",x"00",x"01",x"03", -- 0x0D40
		x"01",x"01",x"00",x"08",x"1D",x"3F",x"3F",x"CE", -- 0x0D48
		x"F7",x"BB",x"F9",x"8F",x"AD",x"71",x"35",x"B6", -- 0x0D50
		x"C4",x"FB",x"FF",x"7D",x"FF",x"F5",x"20",x"10", -- 0x0D58
		x"CC",x"C4",x"66",x"63",x"31",x"39",x"1C",x"1C", -- 0x0D60
		x"04",x"02",x"82",x"C7",x"C3",x"C3",x"E1",x"E0", -- 0x0D68
		x"08",x"08",x"04",x"0E",x"0E",x"87",x"C3",x"E7", -- 0x0D70
		x"63",x"61",x"30",x"38",x"96",x"91",x"C8",x"C8", -- 0x0D78
		x"79",x"0E",x"85",x"80",x"41",x"31",x"0F",x"98", -- 0x0D80
		x"F0",x"FC",x"33",x"00",x"01",x"07",x"8F",x"F7", -- 0x0D88
		x"D8",x"9C",x"9C",x"98",x"0C",x"0E",x"86",x"C7", -- 0x0D90
		x"43",x"20",x"F0",x"78",x"38",x"0C",x"06",x"06", -- 0x0D98
		x"00",x"00",x"C3",x"FF",x"4C",x"04",x"C0",x"E7", -- 0x0DA0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DA8
		x"00",x"E0",x"F0",x"30",x"1C",x"0F",x"C1",x"B8", -- 0x0DB0
		x"CE",x"E3",x"F1",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB8
		x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07", -- 0x0DC0
		x"06",x"0E",x"1C",x"1C",x"3C",x"38",x"78",x"7C", -- 0x0DC8
		x"00",x"01",x"3C",x"6C",x"C8",x"84",x"86",x"42", -- 0x0DD0
		x"43",x"21",x"31",x"30",x"1C",x"1C",x"0E",x"0F", -- 0x0DD8
		x"FE",x"F9",x"F0",x"F0",x"E0",x"F0",x"FD",x"E2", -- 0x0DE0
		x"F2",x"F9",x"D8",x"EC",x"E6",x"F1",x"D0",x"EC", -- 0x0DE8
		x"3F",x"07",x"81",x"C0",x"30",x"0C",x"06",x"E1", -- 0x0DF0
		x"73",x"1E",x"80",x"E0",x"30",x"0C",x"C7",x"70", -- 0x0DF8
		x"E6",x"F3",x"B8",x"E6",x"FB",x"FF",x"FF",x"FF", -- 0x0E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E08
		x"38",x"0F",x"85",x"E0",x"F8",x"FE",x"FF",x"FF", -- 0x0E10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E28
		x"00",x"00",x"01",x"03",x"03",x"03",x"07",x"07", -- 0x0E30
		x"07",x"07",x"0F",x"0F",x"0F",x"1F",x"1F",x"1F", -- 0x0E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0E48
		x"1F",x"1F",x"1F",x"3F",x"3F",x"3F",x"3F",x"7F", -- 0x0E50
		x"7F",x"7F",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x0E58
		x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"BF", -- 0x0E60
		x"4C",x"1C",x"AE",x"1F",x"8F",x"C7",x"FF",x"FF", -- 0x0E68
		x"FF",x"FF",x"7F",x"2F",x"13",x"07",x"AB",x"47", -- 0x0E70
		x"E3",x"73",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E78
		x"FF",x"EF",x"E7",x"E2",x"F1",x"F0",x"FA",x"F4", -- 0x0E80
		x"CE",x"C7",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0E88
		x"FF",x"FF",x"FF",x"FF",x"3F",x"7B",x"B9",x"78", -- 0x0E90
		x"3C",x"1C",x"FE",x"FD",x"F3",x"F1",x"F9",x"FF", -- 0x0E98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"00", -- 0x0EA0
		x"0A",x"80",x"80",x"54",x"EB",x"A8",x"17",x"E5", -- 0x0EA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0EB0
		x"0F",x"40",x"00",x"80",x"60",x"99",x"36",x"6D", -- 0x0EB8
		x"FF",x"FF",x"FF",x"FF",x"17",x"00",x"00",x"40", -- 0x0EC0
		x"F2",x"7D",x"85",x"55",x"6B",x"A8",x"97",x"65", -- 0x0EC8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"01",x"00", -- 0x0ED0
		x"08",x"A0",x"6B",x"96",x"45",x"99",x"36",x"6D", -- 0x0ED8
		x"FF",x"7F",x"01",x"00",x"A6",x"99",x"6C",x"B6", -- 0x0EE0
		x"55",x"AA",x"19",x"B5",x"52",x"49",x"A7",x"9A", -- 0x0EE8
		x"FF",x"FF",x"FF",x"17",x"02",x"00",x"E8",x"E7", -- 0x0EF0
		x"5B",x"B5",x"9F",x"48",x"BA",x"65",x"13",x"96", -- 0x0EF8
		x"00",x"A8",x"4D",x"51",x"26",x"28",x"84",x"B4", -- 0x0F00
		x"05",x"90",x"03",x"CA",x"A8",x"55",x"94",x"65", -- 0x0F08
		x"00",x"00",x"00",x"62",x"98",x"25",x"80",x"9B", -- 0x0F10
		x"25",x"88",x"55",x"28",x"A5",x"52",x"A8",x"13", -- 0x0F18
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F20
		x"FF",x"FF",x"FF",x"3F",x"0F",x"01",x"80",x"44", -- 0x0F28
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F30
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"05", -- 0x0F38
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F40
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F48
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F50
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F60
		x"FF",x"F8",x"C0",x"00",x"00",x"15",x"2A",x"55", -- 0x0F68
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"F8",x"C0", -- 0x0F70
		x"00",x"02",x"06",x"B5",x"0A",x"9A",x"65",x"54", -- 0x0F78
		x"51",x"61",x"B1",x"81",x"21",x"81",x"11",x"A1", -- 0x0F80
		x"51",x"81",x"A1",x"51",x"91",x"61",x"21",x"91", -- 0x0F88
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0F98
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FA0
		x"7F",x"02",x"00",x"00",x"00",x"61",x"BC",x"B6", -- 0x0FA8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0FB0
		x"FF",x"FF",x"37",x"00",x"00",x"00",x"F8",x"A6", -- 0x0FB8
		x"43",x"80",x"00",x"B0",x"52",x"49",x"A7",x"9A", -- 0x0FC0
		x"6A",x"95",x"D2",x"69",x"A6",x"99",x"6C",x"B6", -- 0x0FC8
		x"FF",x"7F",x"1F",x"03",x"00",x"40",x"00",x"94", -- 0x0FD0
		x"68",x"56",x"D1",x"2A",x"D6",x"15",x"E9",x"A6", -- 0x0FD8
		x"A1",x"61",x"81",x"A1",x"61",x"D8",x"90",x"68", -- 0x0FE0
		x"98",x"A6",x"49",x"52",x"B5",x"19",x"AA",x"55", -- 0x0FE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"1F",x"A7", -- 0x0FF0
		x"01",x"00",x"20",x"88",x"40",x"99",x"A5",x"5A", -- 0x0FF8
		x"FF",x"FD",x"FF",x"FF",x"7F",x"BF",x"FF",x"DD", -- 0x1000
		x"F1",x"FB",x"2B",x"EB",x"F7",x"77",x"BF",x"5E", -- 0x1008
		x"FF",x"FF",x"EF",x"DF",x"FD",x"FF",x"FF",x"FF", -- 0x1010
		x"DF",x"DF",x"F7",x"FF",x"FF",x"FF",x"DF",x"FF", -- 0x1018
		x"EE",x"FE",x"F3",x"FF",x"FB",x"EB",x"C9",x"C7", -- 0x1020
		x"85",x"4D",x"5F",x"BF",x"FF",x"5F",x"5D",x"28", -- 0x1028
		x"3F",x"9F",x"9B",x"5F",x"5F",x"7F",x"3D",x"BF", -- 0x1030
		x"FF",x"7F",x"37",x"A3",x"A7",x"AF",x"BF",x"DF", -- 0x1038
		x"6F",x"AB",x"7B",x"7F",x"36",x"7D",x"7B",x"BF", -- 0x1040
		x"DF",x"EF",x"DB",x"D7",x"F6",x"EF",x"ED",x"EF", -- 0x1048
		x"D1",x"D1",x"D3",x"D3",x"D7",x"CF",x"EF",x"ED", -- 0x1050
		x"E9",x"E9",x"EB",x"27",x"37",x"F6",x"F4",x"F4", -- 0x1058
		x"3F",x"BF",x"7F",x"7E",x"BF",x"AF",x"DF",x"EF", -- 0x1060
		x"EB",x"EB",x"F7",x"F7",x"F5",x"FB",x"FF",x"7F", -- 0x1068
		x"FF",x"FF",x"FD",x"FF",x"FF",x"EF",x"F7",x"FF", -- 0x1070
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x1078
		x"7F",x"BE",x"BF",x"BF",x"BF",x"DF",x"D3",x"DF", -- 0x1080
		x"EF",x"EF",x"ED",x"EB",x"F7",x"F5",x"F5",x"F7", -- 0x1088
		x"FF",x"FD",x"9F",x"5F",x"5E",x"7F",x"3F",x"BF", -- 0x1090
		x"67",x"47",x"AF",x"BF",x"DF",x"FF",x"FF",x"FF", -- 0x1098
		x"FE",x"F6",x"E6",x"F9",x"F3",x"FD",x"E2",x"4D", -- 0x10A0
		x"AF",x"FE",x"FF",x"FF",x"DD",x"FD",x"F9",x"F3", -- 0x10A8
		x"7F",x"DF",x"F3",x"E7",x"FF",x"FF",x"7F",x"7F", -- 0x10B0
		x"5B",x"F7",x"F7",x"B7",x"BF",x"AF",x"77",x"EC", -- 0x10B8
		x"FF",x"F7",x"FB",x"BB",x"EE",x"D5",x"EF",x"FA", -- 0x10C0
		x"77",x"BD",x"EB",x"DB",x"FD",x"FE",x"EB",x"F8", -- 0x10C8
		x"F6",x"E7",x"BB",x"7B",x"73",x"FD",x"DD",x"9C", -- 0x10D0
		x"9B",x"6C",x"DF",x"DF",x"7F",x"EF",x"7F",x"B7", -- 0x10D8
		x"4B",x"C7",x"EF",x"DF",x"EF",x"97",x"9F",x"8B", -- 0x10E0
		x"4E",x"A5",x"EF",x"DE",x"FF",x"FF",x"EF",x"FE", -- 0x10E8
		x"DF",x"FF",x"F7",x"FA",x"BA",x"FE",x"9D",x"7E", -- 0x10F0
		x"4F",x"37",x"33",x"9F",x"9A",x"FC",x"BF",x"FF", -- 0x10F8
		x"FF",x"FE",x"F9",x"FF",x"7D",x"BE",x"FE",x"DF", -- 0x1100
		x"DF",x"EF",x"F7",x"F7",x"F7",x"B7",x"3F",x"7F", -- 0x1108
		x"FF",x"EF",x"FF",x"F7",x"F7",x"D7",x"17",x"3F", -- 0x1110
		x"FB",x"7B",x"FB",x"FF",x"BF",x"A7",x"87",x"C7", -- 0x1118
		x"FF",x"FF",x"F7",x"FB",x"BF",x"FF",x"FF",x"FF", -- 0x1120
		x"FF",x"FF",x"FF",x"FF",x"9E",x"8F",x"1F",x"1F", -- 0x1128
		x"FF",x"FF",x"FF",x"BF",x"BF",x"FD",x"FF",x"FF", -- 0x1130
		x"FF",x"FF",x"FF",x"FF",x"0F",x"EF",x"F7",x"FB", -- 0x1138
		x"30",x"60",x"80",x"80",x"C0",x"C0",x"60",x"61", -- 0x1140
		x"37",x"7C",x"83",x"7F",x"FF",x"FF",x"F8",x"E0", -- 0x1148
		x"7F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF", -- 0x1150
		x"1F",x"EF",x"FF",x"F3",x"FF",x"FD",x"7E",x"3F", -- 0x1158
		x"0F",x"98",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1160
		x"E3",x"C6",x"89",x"9F",x"3F",x"7C",x"E0",x"C0", -- 0x1168
		x"FF",x"3F",x"CF",x"F7",x"FB",x"FB",x"FD",x"FE", -- 0x1170
		x"1F",x"EF",x"F7",x"FB",x"9F",x"1D",x"0F",x"0F", -- 0x1178
		x"C0",x"C0",x"63",x"67",x"3F",x"3F",x"1F",x"3F", -- 0x1180
		x"7F",x"FB",x"EF",x"E7",x"C7",x"8F",x"1F",x"1F", -- 0x1188
		x"0F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1190
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F", -- 0x1198
		x"1F",x"23",x"47",x"0F",x"1F",x"3F",x"3F",x"39", -- 0x11A0
		x"73",x"BF",x"3F",x"1C",x"38",x"70",x"E0",x"C0", -- 0x11A8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x11B0
		x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"FF",x"FF", -- 0x11B8
		x"19",x"1F",x"0F",x"07",x"0F",x"0F",x"0F",x"0E", -- 0x11C0
		x"1C",x"1C",x"38",x"20",x"20",x"20",x"40",x"40", -- 0x11C8
		x"FF",x"FF",x"F7",x"E3",x"C1",x"C1",x"E1",x"F3", -- 0x11D0
		x"7F",x"3F",x"3F",x"7F",x"7F",x"FF",x"FF",x"FF", -- 0x11D8
		x"40",x"80",x"81",x"81",x"03",x"03",x"07",x"06", -- 0x11E0
		x"04",x"04",x"04",x"84",x"80",x"89",x"09",x"08", -- 0x11E8
		x"FD",x"F7",x"E3",x"C3",x"C6",x"8F",x"0F",x"0F", -- 0x11F0
		x"0F",x"1D",x"39",x"38",x"36",x"27",x"A1",x"42", -- 0x11F8
		x"FF",x"FF",x"FF",x"FC",x"F8",x"F0",x"E0",x"C0", -- 0x1200
		x"CC",x"86",x"03",x"03",x"06",x"0C",x"0C",x"19", -- 0x1208
		x"C8",x"90",x"31",x"73",x"3E",x"38",x"70",x"64", -- 0x1210
		x"C4",x"C6",x"82",x"01",x"01",x"03",x"C7",x"E7", -- 0x1218
		x"40",x"80",x"80",x"00",x"00",x"00",x"01",x"01", -- 0x1220
		x"00",x"00",x"30",x"19",x"19",x"12",x"10",x"10", -- 0x1228
		x"6F",x"3C",x"38",x"70",x"60",x"E1",x"C3",x"87", -- 0x1230
		x"07",x"87",x"8F",x"0F",x"0F",x"1E",x"1E",x"1C", -- 0x1238
		x"22",x"24",x"24",x"44",x"48",x"48",x"48",x"48", -- 0x1240
		x"88",x"8A",x"84",x"81",x"09",x"08",x"09",x"08", -- 0x1248
		x"1C",x"18",x"38",x"30",x"70",x"E0",x"E0",x"C0", -- 0x1250
		x"80",x"00",x"00",x"00",x"01",x"02",x"02",x"84", -- 0x1258
		x"08",x"08",x"10",x"10",x"00",x"20",x"40",x"40", -- 0x1260
		x"41",x"41",x"80",x"80",x"40",x"40",x"40",x"60", -- 0x1268
		x"24",x"34",x"0C",x"04",x"06",x"08",x"08",x"08", -- 0x1270
		x"08",x"C8",x"70",x"11",x"12",x"22",x"82",x"84", -- 0x1278
		x"01",x"01",x"08",x"06",x"03",x"01",x"21",x"3A", -- 0x1280
		x"1C",x"0C",x"08",x"08",x"08",x"09",x"04",x"04", -- 0x1288
		x"00",x"00",x"B1",x"91",x"11",x"23",x"44",x"24", -- 0x1290
		x"6C",x"9C",x"48",x"48",x"98",x"30",x"90",x"90", -- 0x1298
		x"08",x"08",x"12",x"12",x"24",x"24",x"24",x"24", -- 0x12A0
		x"46",x"42",x"40",x"04",x"24",x"20",x"00",x"12", -- 0x12A8
		x"20",x"40",x"40",x"00",x"00",x"80",x"81",x"81", -- 0x12B0
		x"81",x"01",x"01",x"40",x"40",x"45",x"0F",x"27", -- 0x12B8
		x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x12C0
		x"FF",x"FD",x"FE",x"FF",x"FF",x"BF",x"FF",x"FF", -- 0x12C8
		x"FF",x"BF",x"DF",x"FF",x"FF",x"FB",x"FB",x"FF", -- 0x12D0
		x"FF",x"FF",x"7F",x"FF",x"FE",x"FC",x"F8",x"F0", -- 0x12D8
		x"FF",x"FF",x"FF",x"BF",x"DF",x"FE",x"FC",x"FC", -- 0x12E0
		x"FC",x"F8",x"F8",x"F0",x"F1",x"E0",x"C0",x"80", -- 0x12E8
		x"E0",x"C8",x"C4",x"86",x"03",x"01",x"00",x"01", -- 0x12F0
		x"02",x"42",x"F4",x"3C",x"1C",x"0C",x"08",x"08", -- 0x12F8
		x"C0",x"80",x"90",x"00",x"00",x"03",x"00",x"00", -- 0x1300
		x"00",x"00",x"00",x"00",x"40",x"00",x"00",x"00", -- 0x1308
		x"08",x"10",x"10",x"10",x"30",x"20",x"E0",x"20", -- 0x1310
		x"20",x"40",x"40",x"40",x"40",x"60",x"20",x"30", -- 0x1318
		x"03",x"00",x"00",x"40",x"00",x"00",x"00",x"00", -- 0x1320
		x"04",x"03",x"02",x"02",x"02",x"06",x"02",x"02", -- 0x1328
		x"61",x"C2",x"42",x"4A",x"4E",x"C4",x"84",x"84", -- 0x1330
		x"84",x"04",x"08",x"08",x"08",x"28",x"10",x"10", -- 0x1338
		x"03",x"02",x"02",x"16",x"3C",x"1C",x"0C",x"04", -- 0x1340
		x"04",x"04",x"02",x"02",x"02",x"02",x"32",x"39", -- 0x1348
		x"28",x"78",x"30",x"10",x"50",x"E0",x"20",x"20", -- 0x1350
		x"20",x"20",x"20",x"10",x"10",x"10",x"08",x"08", -- 0x1358
		x"1F",x"0F",x"06",x"22",x"3C",x"0C",x"04",x"04", -- 0x1360
		x"04",x"04",x"02",x"02",x"12",x"1E",x"02",x"00", -- 0x1368
		x"08",x"08",x"04",x"04",x"04",x"08",x"08",x"08", -- 0x1370
		x"08",x"10",x"10",x"D0",x"70",x"10",x"10",x"00", -- 0x1378
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F7",x"FB", -- 0x1380
		x"FF",x"FF",x"FD",x"FE",x"DF",x"FF",x"FF",x"FF", -- 0x1388
		x"FF",x"FF",x"DE",x"FE",x"FC",x"FC",x"FC",x"F8", -- 0x1390
		x"F8",x"F8",x"F8",x"F0",x"F0",x"F0",x"E0",x"E0", -- 0x1398
		x"FF",x"FF",x"FF",x"DF",x"EF",x"FE",x"FF",x"FF", -- 0x13A0
		x"FF",x"FF",x"FF",x"BF",x"FE",x"EE",x"EE",x"FE", -- 0x13A8
		x"C0",x"C0",x"80",x"84",x"80",x"80",x"00",x"00", -- 0x13B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"00", -- 0x13B8
		x"FC",x"FC",x"FC",x"BC",x"DC",x"F8",x"F8",x"F8", -- 0x13C0
		x"F8",x"F8",x"F8",x"B0",x"F0",x"F0",x"F0",x"F0", -- 0x13C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00", -- 0x13D0
		x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00", -- 0x13D8
		x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C4",x"C0", -- 0x13E0
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"E0",x"E0", -- 0x13E8
		x"00",x"00",x"00",x"08",x"04",x"00",x"00",x"00", -- 0x13F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F8
		x"6B",x"AF",x"2E",x"7F",x"57",x"DB",x"7D",x"5C", -- 0x1400
		x"8E",x"7F",x"7F",x"37",x"19",x"78",x"E9",x"29", -- 0x1408
		x"17",x"37",x"37",x"71",x"E0",x"ED",x"EF",x"EF", -- 0x1410
		x"2F",x"63",x"C1",x"D1",x"DB",x"DF",x"DF",x"DF", -- 0x1418
		x"2F",x"47",x"43",x"F3",x"BB",x"7F",x"7D",x"FF", -- 0x1420
		x"FF",x"FB",x"FB",x"FB",x"FF",x"71",x"1A",x"26", -- 0x1428
		x"C6",x"B1",x"BB",x"BF",x"BF",x"3F",x"4F",x"C7", -- 0x1430
		x"AF",x"2D",x"7F",x"7F",x"7F",x"9B",x"9D",x"3F", -- 0x1438
		x"FA",x"B7",x"77",x"F5",x"E9",x"A3",x"DF",x"DF", -- 0x1440
		x"DF",x"BF",x"BF",x"5F",x"8F",x"1F",x"3D",x"7F", -- 0x1448
		x"FF",x"DF",x"FF",x"FF",x"FF",x"F7",x"DF",x"DF", -- 0x1450
		x"FF",x"FF",x"FF",x"FD",x"DF",x"EF",x"FF",x"FF", -- 0x1458
		x"FE",x"FC",x"76",x"77",x"D7",x"1D",x"39",x"3F", -- 0x1460
		x"76",x"66",x"EE",x"FF",x"FF",x"7E",x"7F",x"73", -- 0x1468
		x"FD",x"7E",x"BE",x"BE",x"FF",x"FF",x"4B",x"CB", -- 0x1470
		x"DF",x"FF",x"F7",x"37",x"15",x"3C",x"68",x"F8", -- 0x1478
		x"7F",x"6F",x"F3",x"F7",x"DF",x"FB",x"BF",x"FF", -- 0x1480
		x"FF",x"6F",x"3E",x"5F",x"FD",x"AD",x"DF",x"7A", -- 0x1488
		x"FC",x"FD",x"99",x"B9",x"F3",x"F7",x"FF",x"FF", -- 0x1490
		x"FF",x"FF",x"FF",x"F7",x"FF",x"EF",x"EF",x"7D", -- 0x1498
		x"FF",x"FF",x"BB",x"D1",x"DB",x"FF",x"FF",x"FF", -- 0x14A0
		x"FF",x"FF",x"FD",x"FC",x"F9",x"B9",x"7F",x"FF", -- 0x14A8
		x"F8",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x14B0
		x"FF",x"FF",x"FF",x"FB",x"FB",x"FF",x"FF",x"DF", -- 0x14B8
		x"F4",x"F6",x"FF",x"EF",x"FA",x"D0",x"F2",x"B3", -- 0x14C0
		x"F5",x"FD",x"7F",x"7F",x"35",x"1F",x"AB",x"F3", -- 0x14C8
		x"BB",x"FB",x"7F",x"F7",x"F7",x"FF",x"BF",x"2F", -- 0x14D0
		x"EF",x"FF",x"F9",x"E9",x"FB",x"FF",x"FF",x"D3", -- 0x14D8
		x"F4",x"97",x"B7",x"34",x"3C",x"6D",x"6F",x"6F", -- 0x14E0
		x"7F",x"DF",x"DF",x"FF",x"BF",x"BF",x"BE",x"CF", -- 0x14E8
		x"FF",x"EF",x"A7",x"A3",x"A3",x"B7",x"FF",x"7F", -- 0x14F0
		x"3F",x"AF",x"C7",x"6E",x"6F",x"FF",x"FD",x"7F", -- 0x14F8
		x"4A",x"9A",x"1B",x"1F",x"37",x"37",x"7D",x"6F", -- 0x1500
		x"EF",x"F3",x"F7",x"BF",x"FE",x"4F",x"DF",x"FF", -- 0x1508
		x"7F",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF",x"FF", -- 0x1510
		x"FF",x"F7",x"EF",x"FF",x"FF",x"FD",x"FF",x"FF", -- 0x1518
		x"08",x"08",x"88",x"84",x"B4",x"04",x"04",x"04", -- 0x1520
		x"04",x"06",x"02",x"03",x"81",x"81",x"80",x"C1", -- 0x1528
		x"01",x"00",x"00",x"00",x"20",x"30",x"10",x"18", -- 0x1530
		x"08",x"18",x"2C",x"06",x"03",x"00",x"80",x"80", -- 0x1538
		x"40",x"40",x"20",x"20",x"20",x"30",x"10",x"18", -- 0x1540
		x"08",x"08",x"08",x"0C",x"06",x"0E",x"1F",x"99", -- 0x1548
		x"80",x"80",x"C0",x"40",x"61",x"31",x"1F",x"0F", -- 0x1550
		x"13",x"21",x"00",x"00",x"01",x"00",x"00",x"01", -- 0x1558
		x"80",x"80",x"40",x"20",x"10",x"10",x"88",x"42", -- 0x1560
		x"01",x"20",x"20",x"10",x"08",x"06",x"03",x"01", -- 0x1568
		x"80",x"C1",x"67",x"1D",x"01",x"00",x"00",x"00", -- 0x1570
		x"01",x"83",x"64",x"3E",x"05",x"01",x"07",x"FE", -- 0x1578
		x"10",x"10",x"08",x"04",x"83",x"80",x"C0",x"60", -- 0x1580
		x"30",x"18",x"38",x"3C",x"66",x"E3",x"C0",x"00", -- 0x1588
		x"37",x"07",x"0F",x"1F",x"3F",x"FE",x"7D",x"0B", -- 0x1590
		x"13",x"07",x"0F",x"0F",x"1E",x"BF",x"FF",x"0F", -- 0x1598
		x"00",x"00",x"40",x"20",x"10",x"08",x"06",x"01", -- 0x15A0
		x"00",x"00",x"00",x"00",x"C0",x"60",x"F8",x"EF", -- 0x15A8
		x"0F",x"0F",x"1D",x"13",x"03",x"07",x"0F",x"1D", -- 0x15B0
		x"F3",x"03",x"07",x"0F",x"1F",x"3F",x"3F",x"CB", -- 0x15B8
		x"00",x"00",x"00",x"00",x"00",x"98",x"7C",x"37", -- 0x15C0
		x"21",x"60",x"40",x"40",x"80",x"00",x"00",x"00", -- 0x15C8
		x"77",x"E7",x"0F",x"0F",x"0F",x"1F",x"3F",x"3F", -- 0x15D0
		x"FF",x"3E",x"3E",x"3C",x"30",x"01",x"01",x"00", -- 0x15D8
		x"10",x"18",x"0C",x"06",x"03",x"00",x"00",x"00", -- 0x15E0
		x"00",x"00",x"00",x"00",x"07",x"FF",x"FF",x"FF", -- 0x15E8
		x"03",x"07",x"0F",x"1F",x"FF",x"1B",x"17",x"07", -- 0x15F0
		x"0E",x"1F",x"3F",x"F7",x"EF",x"FF",x"FF",x"FF", -- 0x15F8
		x"12",x"6D",x"A4",x"E4",x"40",x"C6",x"46",x"2F", -- 0x1600
		x"24",x"24",x"24",x"24",x"32",x"11",x"18",x"08", -- 0x1608
		x"61",x"C1",x"40",x"40",x"4F",x"4F",x"87",x"81", -- 0x1610
		x"81",x"81",x"81",x"00",x"C0",x"C0",x"40",x"63", -- 0x1618
		x"1C",x"74",x"48",x"08",x"08",x"08",x"04",x"04", -- 0x1620
		x"06",x"1D",x"39",x"31",x"60",x"C6",x"8F",x"89", -- 0x1628
		x"96",x"94",x"50",x"58",x"48",x"48",x"24",x"24", -- 0x1630
		x"24",x"04",x"16",x"12",x"96",x"85",x"08",x"1C", -- 0x1638
		x"07",x"07",x"06",x"00",x"00",x"00",x"00",x"00", -- 0x1640
		x"00",x"00",x"01",x"01",x"01",x"03",x"02",x"00", -- 0x1648
		x"01",x"00",x"06",x"06",x"04",x"00",x"01",x"03", -- 0x1650
		x"03",x"42",x"E0",x"C0",x"80",x"00",x"08",x"18", -- 0x1658
		x"08",x"09",x"09",x"07",x"8F",x"98",x"98",x"89", -- 0x1660
		x"49",x"49",x"48",x"40",x"44",x"24",x"24",x"22", -- 0x1668
		x"84",x"0E",x"1E",x"3B",x"30",x"00",x"80",x"80", -- 0x1670
		x"80",x"80",x"80",x"40",x"20",x"00",x"10",x"32", -- 0x1678
		x"C2",x"02",x"00",x"00",x"00",x"03",x"07",x"1E", -- 0x1680
		x"1E",x"1C",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1688
		x"63",x"20",x"20",x"00",x"00",x"10",x"10",x"00", -- 0x1690
		x"00",x"0C",x"0C",x"00",x"00",x"00",x"20",x"E0", -- 0x1698
		x"71",x"F8",x"F8",x"7C",x"27",x"01",x"00",x"00", -- 0x16A0
		x"01",x"03",x"03",x"00",x"00",x"20",x"02",x"00", -- 0x16A8
		x"E4",x"C4",x"06",x"03",x"01",x"83",x"87",x"87", -- 0x16B0
		x"C3",x"C3",x"71",x"0C",x"02",x"0D",x"0E",x"06", -- 0x16B8
		x"00",x"80",x"C0",x"C0",x"E0",x"F0",x"F8",x"BC", -- 0x16C0
		x"FE",x"FF",x"FF",x"FF",x"FF",x"DE",x"EF",x"FF", -- 0x16C8
		x"00",x"00",x"40",x"00",x"00",x"00",x"08",x"00", -- 0x16D0
		x"00",x"00",x"C0",x"F0",x"FC",x"FF",x"FF",x"FF", -- 0x16D8
		x"01",x"02",x"02",x"02",x"1A",x"1E",x"3C",x"04", -- 0x16E0
		x"04",x"04",x"04",x"04",x"06",x"02",x"01",x"03", -- 0x16E8
		x"20",x"20",x"E0",x"F1",x"10",x"13",x"13",x"3B", -- 0x16F0
		x"78",x"08",x"08",x"1C",x"24",x"04",x"08",x"38", -- 0x16F8
		x"03",x"02",x"02",x"1A",x"3E",x"3E",x"14",x"04", -- 0x1700
		x"04",x"04",x"04",x"04",x"06",x"02",x"02",x"01", -- 0x1708
		x"38",x"78",x"10",x"70",x"F0",x"20",x"20",x"20", -- 0x1710
		x"20",x"20",x"20",x"10",x"10",x"10",x"08",x"08", -- 0x1718
		x"02",x"02",x"02",x"02",x"02",x"02",x"03",x"00", -- 0x1720
		x"00",x"00",x"01",x"03",x"46",x"00",x"00",x"00", -- 0x1728
		x"70",x"50",x"18",x"18",x"28",x"08",x"04",x"8C", -- 0x1730
		x"8C",x"94",x"C4",x"42",x"46",x"4E",x"4E",x"6F", -- 0x1738
		x"00",x"06",x"07",x"03",x"01",x"00",x"00",x"00", -- 0x1740
		x"00",x"00",x"01",x"03",x"00",x"00",x"00",x"01", -- 0x1748
		x"10",x"20",x"60",x"C3",x"C3",x"46",x"40",x"60", -- 0x1750
		x"20",x"60",x"E0",x"30",x"10",x"10",x"70",x"D8", -- 0x1758
		x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00", -- 0x1760
		x"00",x"00",x"00",x"88",x"80",x"80",x"C0",x"C0", -- 0x1768
		x"C8",x"08",x"0C",x"04",x"04",x"04",x"06",x"02", -- 0x1770
		x"03",x"01",x"03",x"02",x"06",x"04",x"48",x"00", -- 0x1778
		x"C0",x"E0",x"F0",x"F0",x"F8",x"FC",x"BE",x"DE", -- 0x1780
		x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"FF", -- 0x1788
		x"00",x"00",x"00",x"80",x"00",x"00",x"08",x"00", -- 0x1790
		x"00",x"80",x"C0",x"C0",x"E0",x"F8",x"FC",x"FE", -- 0x1798
		x"E0",x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",x"F8", -- 0x17A0
		x"B8",x"F8",x"F8",x"F8",x"FC",x"F4",x"FE",x"FE", -- 0x17A8
		x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00", -- 0x17B0
		x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x17B8
		x"FE",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x17C0
		x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",x"FF",x"FF", -- 0x17C8
		x"00",x"00",x"00",x"00",x"80",x"84",x"80",x"C0", -- 0x17D0
		x"C0",x"C0",x"E0",x"E0",x"E0",x"E0",x"F0",x"F0", -- 0x17D8
		x"FF",x"FF",x"FF",x"FF",x"FB",x"FD",x"FF",x"FF", -- 0x17E0
		x"FF",x"DF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x17E8
		x"F0",x"D8",x"F8",x"FC",x"FC",x"FC",x"FC",x"FC", -- 0x17F0
		x"FE",x"FE",x"FF",x"EF",x"3F",x"FF",x"FF",x"FF", -- 0x17F8
		x"FF",x"FE",x"FF",x"F7",x"F7",x"FE",x"FF",x"FF", -- 0x1800
		x"FF",x"FF",x"FF",x"DF",x"FF",x"FF",x"FE",x"FF", -- 0x1808
		x"91",x"25",x"72",x"DA",x"5C",x"2E",x"9F",x"4C", -- 0x1810
		x"AE",x"DA",x"76",x"83",x"E5",x"A2",x"D1",x"F0", -- 0x1818
		x"95",x"12",x"4A",x"2E",x"59",x"DC",x"26",x"66", -- 0x1820
		x"0B",x"41",x"87",x"E1",x"D5",x"F5",x"BA",x"FF", -- 0x1828
		x"81",x"A5",x"F2",x"D2",x"54",x"2E",x"5F",x"CC", -- 0x1830
		x"6E",x"DA",x"B7",x"83",x"05",x"42",x"D1",x"F0", -- 0x1838
		x"9D",x"2E",x"04",x"84",x"42",x"D4",x"FA",x"D8", -- 0x1840
		x"E1",x"E4",x"C3",x"E9",x"F3",x"FD",x"B2",x"FE", -- 0x1848
		x"81",x"A5",x"D2",x"52",x"14",x"6E",x"3F",x"CC", -- 0x1850
		x"5E",x"DA",x"F6",x"C0",x"5A",x"5F",x"DF",x"0A", -- 0x1858
		x"95",x"12",x"4A",x"2E",x"99",x"9F",x"A6",x"66", -- 0x1860
		x"0B",x"A0",x"D7",x"E0",x"EC",x"FA",x"FF",x"FE", -- 0x1868
		x"81",x"A5",x"D2",x"D3",x"15",x"6E",x"1F",x"AD", -- 0x1870
		x"6F",x"DA",x"B6",x"C2",x"47",x"E3",x"D1",x"FC", -- 0x1878
		x"95",x"12",x"4A",x"86",x"4B",x"D2",x"90",x"EC", -- 0x1880
		x"F9",x"FE",x"BD",x"FF",x"FF",x"FF",x"F6",x"FF", -- 0x1888
		x"81",x"A5",x"D2",x"D2",x"14",x"6E",x"3F",x"8C", -- 0x1890
		x"2C",x"D5",x"2B",x"9F",x"FD",x"FF",x"EF",x"FF", -- 0x1898
		x"95",x"13",x"4B",x"2F",x"9F",x"9F",x"27",x"67", -- 0x18A0
		x"0B",x"E7",x"FF",x"4F",x"BD",x"1F",x"3F",x"7F", -- 0x18A8
		x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD", -- 0x18B0
		x"FF",x"BF",x"FF",x"FF",x"EF",x"FB",x"FB",x"DF", -- 0x18B8
		x"7C",x"DB",x"B9",x"12",x"01",x"47",x"CB",x"59", -- 0x18C0
		x"4F",x"73",x"B9",x"7A",x"BA",x"57",x"B7",x"3F", -- 0x18C8
		x"74",x"BA",x"D7",x"EF",x"6F",x"5E",x"AB",x"D2", -- 0x18D0
		x"85",x"57",x"6F",x"7F",x"FF",x"FF",x"FF",x"FF", -- 0x18D8
		x"95",x"12",x"4A",x"2E",x"98",x"9F",x"26",x"66", -- 0x18E0
		x"0B",x"A1",x"F7",x"69",x"BB",x"25",x"71",x"5B", -- 0x18E8
		x"81",x"A7",x"D3",x"DB",x"17",x"6F",x"BF",x"CF", -- 0x18F0
		x"57",x"EF",x"8D",x"FF",x"7F",x"7F",x"7B",x"FF", -- 0x18F8
		x"95",x"12",x"4A",x"2C",x"9C",x"9E",x"27",x"66", -- 0x1900
		x"0A",x"AF",x"FF",x"4D",x"BF",x"1F",x"3F",x"7F", -- 0x1908
		x"81",x"A5",x"D3",x"D3",x"15",x"67",x"37",x"7D", -- 0x1910
		x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"FF", -- 0x1918
		x"95",x"12",x"4A",x"2C",x"8A",x"9F",x"36",x"72", -- 0x1920
		x"3B",x"FF",x"BF",x"FF",x"FF",x"FF",x"EF",x"FF", -- 0x1928
		x"81",x"A5",x"D3",x"D3",x"15",x"67",x"37",x"BF", -- 0x1930
		x"FF",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1938
		x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1940
		x"DF",x"FF",x"FF",x"FF",x"FE",x"FD",x"FE",x"FE", -- 0x1948
		x"FA",x"EE",x"C7",x"FB",x"9D",x"E7",x"C6",x"B2", -- 0x1950
		x"E0",x"D0",x"69",x"95",x"55",x"78",x"94",x"32", -- 0x1958
		x"FF",x"FF",x"FF",x"FF",x"F1",x"FF",x"EB",x"D9", -- 0x1960
		x"4F",x"73",x"BD",x"7B",x"B2",x"5C",x"CA",x"64", -- 0x1968
		x"FF",x"FE",x"FB",x"9F",x"4F",x"5E",x"AB",x"D2", -- 0x1970
		x"84",x"70",x"7C",x"2E",x"3F",x"4E",x"36",x"0C", -- 0x1978
		x"FF",x"FF",x"F8",x"FE",x"F5",x"FD",x"E3",x"E9", -- 0x1980
		x"F3",x"EB",x"D1",x"DB",x"B2",x"BD",x"2A",x"04", -- 0x1988
		x"74",x"9A",x"D7",x"CF",x"6F",x"5E",x"AB",x"D2", -- 0x1990
		x"84",x"60",x"64",x"2E",x"3F",x"4E",x"36",x"0C", -- 0x1998
		x"FF",x"DF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF", -- 0x19A0
		x"FF",x"FB",x"FD",x"FD",x"BA",x"D5",x"CA",x"64", -- 0x19A8
		x"FC",x"F8",x"F9",x"FF",x"BF",x"9E",x"4B",x"B2", -- 0x19B0
		x"84",x"70",x"7C",x"2E",x"3F",x"4E",x"36",x"0C", -- 0x19B8
		x"FF",x"FF",x"BF",x"FF",x"FF",x"FB",x"FF",x"FF", -- 0x19C0
		x"FF",x"FE",x"FF",x"FD",x"FE",x"EC",x"4A",x"67", -- 0x19C8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF", -- 0x19D0
		x"F8",x"F2",x"6A",x"16",x"15",x"78",x"94",x"32", -- 0x19D8
		x"AF",x"7F",x"B7",x"6B",x"B3",x"55",x"FE",x"18", -- 0x19E0
		x"4F",x"73",x"B1",x"7A",x"B1",x"5E",x"CB",x"67", -- 0x19E8
		x"FF",x"FF",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x19F0
		x"FF",x"FF",x"F7",x"F7",x"7F",x"FF",x"FF",x"FF", -- 0x19F8
		x"FF",x"7F",x"BF",x"7B",x"B1",x"57",x"FB",x"59", -- 0x1A00
		x"4F",x"73",x"B9",x"7B",x"B2",x"5C",x"CA",x"67", -- 0x1A08
		x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"FF",x"FF", -- 0x1A10
		x"BF",x"53",x"2B",x"96",x"D5",x"78",x"94",x"32", -- 0x1A18
		x"49",x"2B",x"BF",x"7A",x"B1",x"57",x"FB",x"59", -- 0x1A20
		x"4F",x"73",x"B9",x"7B",x"B3",x"5D",x"CA",x"67", -- 0x1A28
		x"FF",x"FF",x"FF",x"7F",x"7F",x"7F",x"FF",x"FF", -- 0x1A30
		x"A7",x"63",x"2F",x"17",x"97",x"FF",x"97",x"33", -- 0x1A38
		x"EF",x"7F",x"BF",x"6B",x"B3",x"55",x"FB",x"19", -- 0x1A40
		x"4F",x"73",x"B1",x"7B",x"B0",x"5E",x"CA",x"67", -- 0x1A48
		x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1A50
		x"FF",x"FF",x"FF",x"5F",x"17",x"79",x"95",x"32", -- 0x1A58
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"B9", -- 0x1A60
		x"6F",x"53",x"B9",x"6F",x"B2",x"58",x"CA",x"67", -- 0x1A68
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F", -- 0x1A70
		x"FF",x"DF",x"5F",x"97",x"17",x"7F",x"97",x"33", -- 0x1A78
		x"FF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7", -- 0x1A80
		x"CB",x"A1",x"F7",x"71",x"BB",x"25",x"71",x"5B", -- 0x1A88
		x"FF",x"FF",x"FF",x"FF",x"F7",x"FF",x"FF",x"EF", -- 0x1A90
		x"5E",x"DB",x"F7",x"C1",x"4A",x"6F",x"FF",x"4A", -- 0x1A98
		x"95",x"12",x"4B",x"2E",x"9B",x"9D",x"20",x"74", -- 0x1AA0
		x"3D",x"FF",x"FE",x"FB",x"FF",x"FF",x"FF",x"FF", -- 0x1AA8
		x"81",x"25",x"D2",x"DA",x"1C",x"6E",x"BF",x"1C", -- 0x1AB0
		x"1E",x"9A",x"75",x"97",x"FF",x"F7",x"FF",x"FF", -- 0x1AB8
		x"FE",x"FC",x"FE",x"FD",x"F8",x"FC",x"BE",x"FE", -- 0x1AC0
		x"FD",x"F8",x"FF",x"FC",x"FD",x"F8",x"FC",x"FE", -- 0x1AC8
		x"81",x"25",x"52",x"DA",x"1C",x"6E",x"3F",x"CC", -- 0x1AD0
		x"5E",x"DA",x"F6",x"D0",x"6A",x"57",x"DF",x"0A", -- 0x1AD8
		x"4B",x"2D",x"B9",x"7A",x"B1",x"57",x"FB",x"59", -- 0x1AE0
		x"4F",x"73",x"B9",x"7A",x"B3",x"5D",x"CB",x"67", -- 0x1AE8
		x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FB", -- 0x1AF0
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1AF8
		x"BF",x"BB",x"FF",x"FA",x"DF",x"FF",x"FB",x"EF", -- 0x1B00
		x"EF",x"EF",x"FF",x"BF",x"BB",x"BB",x"FF",x"FF", -- 0x1B08
		x"7D",x"75",x"FF",x"DB",x"DB",x"7B",x"7F",x"DD", -- 0x1B10
		x"DD",x"7F",x"EF",x"EF",x"FF",x"FB",x"7B",x"7E", -- 0x1B18
		x"FF",x"FB",x"BB",x"FF",x"FF",x"FE",x"DC",x"DD", -- 0x1B20
		x"FD",x"FF",x"EF",x"ED",x"FF",x"FF",x"F7",x"FF", -- 0x1B28
		x"7F",x"FB",x"FB",x"DB",x"FF",x"FF",x"FF",x"DF", -- 0x1B30
		x"DF",x"F7",x"FF",x"FE",x"7E",x"7F",x"EF",x"EF", -- 0x1B38
		x"FF",x"FB",x"BB",x"FF",x"FF",x"FE",x"DC",x"DD", -- 0x1B40
		x"FD",x"FF",x"EF",x"ED",x"FF",x"FF",x"F7",x"FF", -- 0x1B48
		x"7C",x"FA",x"FB",x"DA",x"FF",x"FF",x"FF",x"DF", -- 0x1B50
		x"DF",x"F7",x"FF",x"FE",x"7E",x"7F",x"EF",x"EF", -- 0x1B58
		x"7C",x"DB",x"B9",x"13",x"41",x"27",x"8B",x"59", -- 0x1B60
		x"4F",x"73",x"B1",x"7B",x"B2",x"5C",x"CA",x"64", -- 0x1B68
		x"74",x"BA",x"D7",x"DF",x"4F",x"5E",x"AB",x"D2", -- 0x1B70
		x"84",x"60",x"64",x"2E",x"3F",x"4E",x"36",x"0C", -- 0x1B78
		x"95",x"12",x"4A",x"2E",x"99",x"9C",x"26",x"66", -- 0x1B80
		x"0B",x"A1",x"F7",x"61",x"B3",x"25",x"71",x"5B", -- 0x1B88
		x"81",x"A5",x"D2",x"D2",x"14",x"6E",x"3F",x"CC", -- 0x1B90
		x"5E",x"DA",x"F6",x"C0",x"5A",x"5F",x"DF",x"0A", -- 0x1B98
		x"49",x"2D",x"BC",x"7A",x"B1",x"57",x"FB",x"59", -- 0x1BA0
		x"4F",x"73",x"B1",x"7B",x"B2",x"5C",x"CA",x"67", -- 0x1BA8
		x"A6",x"EF",x"DF",x"5B",x"5D",x"4F",x"A4",x"C0", -- 0x1BB0
		x"84",x"66",x"2A",x"16",x"15",x"78",x"94",x"32", -- 0x1BB8
		x"FF",x"FF",x"FF",x"FF",x"EF",x"E7",x"E2",x"F1", -- 0x1BC0
		x"F0",x"FA",x"F4",x"CE",x"C7",x"E7",x"FF",x"FF", -- 0x1BC8
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"38", -- 0x1BD0
		x"78",x"B8",x"78",x"38",x"18",x"F8",x"F8",x"F8", -- 0x1BD8
		x"FF",x"FF",x"FF",x"FF",x"EF",x"E7",x"E2",x"F1", -- 0x1BE0
		x"F0",x"FA",x"F4",x"CE",x"C7",x"E7",x"FF",x"FF", -- 0x1BE8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F", -- 0x1BF0
		x"7F",x"BF",x"7F",x"3F",x"1F",x"FF",x"FF",x"FF", -- 0x1BF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"1F", -- 0x1C08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"01",x"FD", -- 0x1C18
		x"FF",x"FF",x"4A",x"73",x"00",x"00",x"F3",x"08", -- 0x1C20
		x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C", -- 0x1C28
		x"F8",x"00",x"53",x"9F",x"01",x"00",x"FC",x"07", -- 0x1C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C38
		x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C", -- 0x1C40
		x"0C",x"FF",x"00",x"00",x"3E",x"00",x"00",x"00", -- 0x1C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C50
		x"03",x"FC",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1C58
		x"00",x"00",x"00",x"00",x"00",x"2F",x"E0",x"1F", -- 0x1C60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C68
		x"00",x"20",x"40",x"00",x"00",x"BE",x"00",x"FF", -- 0x1C70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C78
		x"FF",x"FE",x"8E",x"BC",x"5C",x"3F",x"9F",x"7F", -- 0x1C80
		x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C88
		x"0F",x"27",x"5F",x"AF",x"FF",x"FF",x"FF",x"FF", -- 0x1C90
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1C98
		x"FF",x"07",x"01",x"FD",x"7D",x"7D",x"61",x"00", -- 0x1CA0
		x"0F",x"1F",x"3F",x"3F",x"3E",x"3E",x"3E",x"27", -- 0x1CA8
		x"F9",x"FF",x"FF",x"FF",x"FF",x"80",x"3F",x"7F", -- 0x1CB0
		x"F8",x"E3",x"0C",x"18",x"10",x"80",x"00",x"C0", -- 0x1CB8
		x"04",x"04",x"01",x"00",x"00",x"00",x"00",x"10", -- 0x1CC0
		x"08",x"04",x"02",x"01",x"00",x"00",x"80",x"40", -- 0x1CC8
		x"50",x"10",x"10",x"50",x"10",x"10",x"18",x"08", -- 0x1CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1CD8
		x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"7D", -- 0x1CE0
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F7", -- 0x1CF0
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1CF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"81",x"FE", -- 0x1D08
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x1D10
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8", -- 0x1D18
		x"FE",x"E0",x"CF",x"8F",x"08",x"08",x"08",x"03", -- 0x1D20
		x"1C",x"40",x"80",x"00",x"00",x"00",x"00",x"00", -- 0x1D28
		x"FF",x"00",x"FF",x"FF",x"FF",x"E0",x"1F",x"F0", -- 0x1D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D38
		x"00",x"00",x"00",x"00",x"00",x"80",x"E0",x"3E", -- 0x1D40
		x"03",x"00",x"00",x"07",x"00",x"00",x"00",x"00", -- 0x1D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1D50
		x"C0",x"3F",x"00",x"80",x"00",x"00",x"00",x"00", -- 0x1D58
		x"C0",x"00",x"00",x"00",x"00",x"00",x"EF",x"00", -- 0x1D60
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D68
		x"00",x"00",x"2A",x"00",x"00",x"00",x"BE",x"00", -- 0x1D70
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D78
		x"A5",x"F0",x"E2",x"E5",x"CA",x"CF",x"FF",x"FF", -- 0x1D80
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D88
		x"7F",x"FF",x"73",x"E7",x"E3",x"E9",x"FC",x"F8", -- 0x1D90
		x"F9",x"F2",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1D98
		x"FC",x"F0",x"E0",x"E0",x"C0",x"C0",x"C0",x"C0", -- 0x1DA0
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x1DA8
		x"1F",x"20",x"00",x"03",x"00",x"04",x"03",x"00", -- 0x1DB0
		x"00",x"00",x"1E",x"0E",x"00",x"00",x"00",x"00", -- 0x1DB8
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x1DC0
		x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x1DC8
		x"3C",x"3C",x"30",x"3C",x"3C",x"3C",x"3C",x"38", -- 0x1DD0
		x"38",x"38",x"20",x"04",x"08",x"00",x"02",x"00", -- 0x1DD8
		x"E0",x"F0",x"F0",x"F8",x"F8",x"FC",x"FE",x"00", -- 0x1DE0
		x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1DF0
		x"7F",x"80",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1DF8
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E00
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"FF", -- 0x1E08
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1E10
		x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"01",x"FD", -- 0x1E18
		x"FF",x"C0",x"C0",x"C0",x"C0",x"E0",x"00",x"E0", -- 0x1E20
		x"F8",x"00",x"00",x"0F",x"3E",x"7C",x"7C",x"72", -- 0x1E28
		x"FD",x"1F",x"1F",x"15",x"0C",x"0F",x"06",x"00", -- 0x1E30
		x"00",x"70",x"C0",x"01",x"83",x"82",x"82",x"02", -- 0x1E38
		x"72",x"72",x"72",x"72",x"70",x"3E",x"1E",x"06", -- 0x1E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E48
		x"00",x"02",x"02",x"03",x"01",x"00",x"00",x"00", -- 0x1E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1E58
		x"FF",x"BF",x"DF",x"DF",x"FF",x"AB",x"CF",x"8B", -- 0x1E60
		x"32",x"D6",x"65",x"5D",x"37",x"75",x"55",x"DF", -- 0x1E68
		x"FF",x"75",x"7B",x"FF",x"D7",x"CE",x"59",x"29", -- 0x1E70
		x"14",x"61",x"AB",x"7E",x"95",x"DD",x"5B",x"FB", -- 0x1E78
		x"63",x"27",x"8B",x"62",x"DA",x"A6",x"76",x"49", -- 0x1E80
		x"6F",x"AA",x"B9",x"AD",x"A7",x"ED",x"7D",x"7E", -- 0x1E88
		x"FF",x"75",x"FB",x"AF",x"9D",x"17",x"D5",x"A3", -- 0x1E90
		x"68",x"95",x"6D",x"6B",x"6E",x"F6",x"D4",x"DF", -- 0x1E98
		x"EE",x"7A",x"72",x"5D",x"D7",x"DE",x"BB",x"BB", -- 0x1EA0
		x"AB",x"E6",x"D7",x"D5",x"D5",x"7D",x"6F",x"6F", -- 0x1EA8
		x"7F",x"95",x"A3",x"93",x"36",x"CC",x"24",x"DD", -- 0x1EB0
		x"6A",x"5D",x"59",x"AF",x"BD",x"B5",x"D5",x"D7", -- 0x1EB8
		x"7A",x"69",x"EE",x"AB",x"BF",x"2A",x"7F",x"B5", -- 0x1EC0
		x"B7",x"F5",x"FD",x"CC",x"6E",x"6E",x"77",x"75", -- 0x1EC8
		x"7F",x"37",x"47",x"8D",x"4A",x"DE",x"AB",x"57", -- 0x1ED0
		x"DD",x"6B",x"C3",x"B7",x"D3",x"2F",x"83",x"BD", -- 0x1ED8
		x"7F",x"2F",x"AB",x"66",x"42",x"6A",x"51",x"A0", -- 0x1EE0
		x"9B",x"57",x"59",x"52",x"DD",x"B4",x"95",x"DD", -- 0x1EE8
		x"FF",x"75",x"FB",x"7F",x"BD",x"7F",x"F7",x"53", -- 0x1EF0
		x"C5",x"2F",x"A7",x"57",x"E9",x"BF",x"51",x"6D", -- 0x1EF8
		x"FF",x"BF",x"DF",x"DF",x"FF",x"BB",x"6F",x"7F", -- 0x1F00
		x"67",x"96",x"44",x"A9",x"82",x"A0",x"54",x"6E", -- 0x1F08
		x"FF",x"75",x"7B",x"BF",x"9D",x"DF",x"FF",x"FB", -- 0x1F10
		x"FD",x"DF",x"BF",x"37",x"5D",x"B7",x"EF",x"9F", -- 0x1F18
		x"7F",x"37",x"27",x"29",x"D7",x"07",x"BC",x"81", -- 0x1F20
		x"C6",x"A9",x"BC",x"43",x"52",x"EC",x"B2",x"D0", -- 0x1F28
		x"FD",x"7F",x"B5",x"3B",x"FB",x"FD",x"DF",x"FF", -- 0x1F30
		x"EF",x"FF",x"FF",x"BD",x"FB",x"FD",x"7F",x"36", -- 0x1F38
		x"D6",x"BC",x"6E",x"5D",x"95",x"BE",x"E9",x"DA", -- 0x1F40
		x"B2",x"BD",x"5E",x"F7",x"DE",x"7A",x"FE",x"BA", -- 0x1F48
		x"76",x"3F",x"BD",x"9B",x"3D",x"FF",x"3F",x"EF", -- 0x1F50
		x"FF",x"5F",x"3D",x"3B",x"1B",x"95",x"3F",x"7D", -- 0x1F58
		x"FF",x"BF",x"FF",x"FB",x"B9",x"54",x"CF",x"57", -- 0x1F60
		x"09",x"D6",x"A4",x"D6",x"7A",x"7F",x"B6",x"B6", -- 0x1F68
		x"FF",x"B7",x"FF",x"EF",x"FD",x"F7",x"F7",x"DB", -- 0x1F70
		x"EF",x"4B",x"A6",x"2B",x"DB",x"66",x"FD",x"DD", -- 0x1F78
		x"D6",x"96",x"4D",x"EB",x"9F",x"75",x"C6",x"56", -- 0x1F80
		x"3A",x"E0",x"AE",x"FC",x"D5",x"4A",x"A7",x"C6", -- 0x1F88
		x"5C",x"AA",x"EF",x"55",x"5E",x"4A",x"8F",x"AD", -- 0x1F90
		x"B6",x"D6",x"5F",x"CD",x"AF",x"E2",x"AB",x"99", -- 0x1F98
		x"99",x"D5",x"47",x"F5",x"B3",x"FA",x"6A",x"4D", -- 0x1FA0
		x"B5",x"51",x"50",x"5A",x"6A",x"2E",x"35",x"D6", -- 0x1FA8
		x"03",x"C5",x"52",x"AA",x"3E",x"55",x"07",x"5C", -- 0x1FB0
		x"6A",x"60",x"AE",x"F9",x"57",x"32",x"69",x"6B", -- 0x1FB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BE", -- 0x1FC0
		x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"7B",x"80", -- 0x1FD0
		x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FD8
		x"E7",x"CF",x"C6",x"D2",x"F8",x"F1",x"F2",x"E5", -- 0x1FE0
		x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x1FE8
		x"F8",x"18",x"78",x"B8",x"78",x"38",x"F8",x"78", -- 0x1FF0
		x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8"  -- 0x1FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
