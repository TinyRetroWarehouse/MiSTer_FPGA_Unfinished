-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

entity ROM_M7 is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_M7 is


	type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"DC",x"98",x"BA",x"85",x"C0",x"88",x"DC",x"98", -- 0x0000
		x"C8",x"8D",x"CE",x"90",x"D4",x"93",x"DA",x"96", -- 0x0008
		x"DC",x"98",x"36",x"83",x"3C",x"86",x"DC",x"98", -- 0x0010
		x"44",x"8B",x"4A",x"8E",x"50",x"91",x"56",x"94", -- 0x0018
		x"34",x"81",x"B8",x"83",x"BE",x"86",x"42",x"89", -- 0x0020
		x"C6",x"8B",x"CC",x"8E",x"D2",x"91",x"D8",x"94", -- 0x0028
		x"00",x"00",x"65",x"02",x"66",x"02",x"00",x"00", -- 0x0030
		x"01",x"00",x"39",x"02",x"3A",x"02",x"71",x"42", -- 0x0038
		x"02",x"00",x"3B",x"02",x"3C",x"02",x"67",x"02", -- 0x0040
		x"03",x"00",x"3D",x"02",x"3E",x"02",x"68",x"02", -- 0x0048
		x"00",x"00",x"3F",x"02",x"40",x"02",x"69",x"02", -- 0x0050
		x"01",x"00",x"41",x"02",x"42",x"02",x"6A",x"02", -- 0x0058
		x"02",x"00",x"43",x"02",x"44",x"02",x"6B",x"02", -- 0x0060
		x"03",x"00",x"45",x"02",x"46",x"02",x"6C",x"02", -- 0x0068
		x"00",x"00",x"47",x"02",x"48",x"02",x"6D",x"02", -- 0x0070
		x"01",x"00",x"49",x"02",x"4A",x"02",x"4B",x"02", -- 0x0078
		x"02",x"00",x"4C",x"02",x"4D",x"02",x"4E",x"02", -- 0x0080
		x"03",x"00",x"4F",x"02",x"50",x"02",x"51",x"02", -- 0x0088
		x"00",x"00",x"52",x"02",x"53",x"02",x"54",x"02", -- 0x0090
		x"01",x"00",x"55",x"02",x"56",x"02",x"6F",x"02", -- 0x0098
		x"02",x"00",x"57",x"02",x"58",x"02",x"70",x"02", -- 0x00A0
		x"03",x"00",x"59",x"02",x"5A",x"02",x"6E",x"02", -- 0x00A8
		x"FF",x"FF",x"00",x"00",x"5B",x"02",x"5C",x"02", -- 0x00B0
		x"71",x"02",x"01",x"00",x"5D",x"02",x"5E",x"02", -- 0x00B8
		x"03",x"00",x"02",x"00",x"5F",x"02",x"60",x"02", -- 0x00C0
		x"00",x"00",x"03",x"00",x"61",x"02",x"62",x"02", -- 0x00C8
		x"01",x"00",x"00",x"00",x"63",x"02",x"64",x"02", -- 0x00D0
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x00D8
		x"03",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x00E0
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x00E8
		x"01",x"00",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x00F0
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x00F8
		x"03",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x0100
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x0108
		x"01",x"00",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x0110
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x0118
		x"03",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x0120
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x0128
		x"01",x"00",x"FF",x"FF",x"00",x"00",x"03",x"00", -- 0x0130
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0138
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0140
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0148
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0150
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0158
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0160
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0168
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0170
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0178
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0180
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0188
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0190
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0198
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x01A0
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x01A8
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x01B0
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x01B8
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x01C0
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x01C8
		x"02",x"00",x"01",x"00",x"04",x"00",x"05",x"00", -- 0x01D0
		x"01",x"00",x"02",x"00",x"06",x"00",x"07",x"00", -- 0x01D8
		x"00",x"00",x"03",x"00",x"08",x"00",x"09",x"00", -- 0x01E0
		x"03",x"00",x"00",x"00",x"0A",x"00",x"0B",x"00", -- 0x01E8
		x"02",x"00",x"01",x"00",x"0C",x"00",x"0D",x"00", -- 0x01F0
		x"0E",x"00",x"02",x"00",x"72",x"02",x"10",x"00", -- 0x01F8
		x"11",x"00",x"03",x"00",x"12",x"00",x"13",x"00", -- 0x0200
		x"14",x"00",x"00",x"00",x"15",x"00",x"16",x"00", -- 0x0208
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0210
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0218
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0220
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0228
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0230
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0238
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0240
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0248
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0250
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0258
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0260
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0268
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0270
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0278
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0280
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0288
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0290
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0298
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x02A0
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x02A8
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x02B0
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x02B8
		x"14",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x02C0
		x"17",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x02C8
		x"02",x"00",x"0E",x"00",x"00",x"00",x"03",x"00", -- 0x02D0
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x02D8
		x"00",x"00",x"11",x"00",x"02",x"00",x"01",x"00", -- 0x02E0
		x"18",x"00",x"19",x"00",x"03",x"00",x"00",x"00", -- 0x02E8
		x"1A",x"00",x"20",x"00",x"00",x"00",x"03",x"00", -- 0x02F0
		x"1B",x"00",x"21",x"00",x"01",x"00",x"02",x"00", -- 0x02F8
		x"1C",x"00",x"22",x"00",x"02",x"00",x"01",x"00", -- 0x0300
		x"1D",x"00",x"1E",x"00",x"03",x"00",x"00",x"00", -- 0x0308
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0310
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0318
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0320
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0328
		x"02",x"00",x"01",x"00",x"FF",x"FF",x"00",x"00", -- 0x0330
		x"03",x"00",x"01",x"00",x"02",x"00",x"01",x"00", -- 0x0338
		x"02",x"00",x"00",x"00",x"03",x"00",x"02",x"00", -- 0x0340
		x"01",x"00",x"03",x"00",x"00",x"00",x"03",x"00", -- 0x0348
		x"00",x"00",x"02",x"00",x"01",x"00",x"00",x"00", -- 0x0350
		x"03",x"00",x"01",x"00",x"02",x"00",x"01",x"00", -- 0x0358
		x"24",x"00",x"00",x"00",x"03",x"00",x"25",x"00", -- 0x0360
		x"26",x"00",x"27",x"00",x"00",x"00",x"28",x"00", -- 0x0368
		x"6D",x"00",x"29",x"00",x"01",x"00",x"2A",x"00", -- 0x0370
		x"2A",x"80",x"2C",x"00",x"2D",x"00",x"2E",x"00", -- 0x0378
		x"2F",x"00",x"2A",x"00",x"30",x"00",x"70",x"00", -- 0x0380
		x"31",x"00",x"32",x"00",x"2B",x"00",x"71",x"00", -- 0x0388
		x"72",x"00",x"33",x"00",x"74",x"00",x"73",x"00", -- 0x0390
		x"70",x"00",x"34",x"00",x"75",x"00",x"36",x"00", -- 0x0398
		x"37",x"00",x"35",x"00",x"76",x"00",x"38",x"00", -- 0x03A0
		x"39",x"00",x"77",x"00",x"74",x"00",x"75",x"00", -- 0x03A8
		x"76",x"00",x"74",x"00",x"77",x"00",x"FF",x"FF", -- 0x03B0
		x"74",x"00",x"75",x"00",x"76",x"00",x"77",x"00", -- 0x03B8
		x"77",x"00",x"76",x"00",x"75",x"00",x"74",x"00", -- 0x03C0
		x"75",x"00",x"3A",x"00",x"3B",x"00",x"75",x"00", -- 0x03C8
		x"3C",x"00",x"3D",x"00",x"3E",x"00",x"76",x"00", -- 0x03D0
		x"3F",x"00",x"71",x"00",x"40",x"00",x"77",x"00", -- 0x03D8
		x"41",x"00",x"42",x"00",x"43",x"00",x"74",x"00", -- 0x03E0
		x"44",x"00",x"45",x"00",x"46",x"00",x"47",x"00", -- 0x03E8
		x"2D",x"02",x"2D",x"02",x"48",x"00",x"4B",x"00", -- 0x03F0
		x"2D",x"02",x"2D",x"02",x"49",x"00",x"4A",x"00", -- 0x03F8
		x"2D",x"02",x"4C",x"00",x"33",x"00",x"75",x"00", -- 0x0400
		x"4D",x"00",x"4E",x"00",x"34",x"00",x"76",x"00", -- 0x0408
		x"36",x"00",x"37",x"00",x"35",x"00",x"77",x"00", -- 0x0410
		x"38",x"00",x"39",x"00",x"74",x"00",x"75",x"00", -- 0x0418
		x"76",x"00",x"77",x"00",x"75",x"00",x"74",x"00", -- 0x0420
		x"75",x"00",x"76",x"00",x"77",x"00",x"76",x"00", -- 0x0428
		x"74",x"00",x"75",x"00",x"76",x"00",x"77",x"00", -- 0x0430
		x"74",x"00",x"75",x"00",x"3C",x"00",x"3B",x"00", -- 0x0438
		x"76",x"00",x"77",x"00",x"4F",x"00",x"3E",x"00", -- 0x0440
		x"75",x"00",x"3C",x"00",x"3D",x"00",x"72",x"00", -- 0x0448
		x"3C",x"00",x"3F",x"00",x"73",x"00",x"70",x"00", -- 0x0450
		x"3F",x"00",x"50",x"00",x"51",x"00",x"71",x"00", -- 0x0458
		x"52",x"00",x"2D",x"02",x"53",x"00",x"72",x"00", -- 0x0460
		x"54",x"00",x"44",x"40",x"51",x"40",x"55",x"00", -- 0x0468
		x"54",x"40",x"56",x"00",x"57",x"00",x"2D",x"02", -- 0x0470
		x"52",x"40",x"59",x"C0",x"53",x"80",x"2D",x"02", -- 0x0478
		x"73",x"00",x"55",x"40",x"58",x"00",x"2D",x"02", -- 0x0480
		x"5A",x"00",x"37",x"00",x"59",x"00",x"2D",x"02", -- 0x0488
		x"74",x"00",x"5B",x"00",x"59",x"40",x"2D",x"02", -- 0x0490
		x"75",x"00",x"5C",x"00",x"5D",x"00",x"5D",x"80", -- 0x0498
		x"76",x"00",x"5E",x"00",x"5F",x"00",x"5F",x"80", -- 0x04A0
		x"77",x"00",x"74",x"00",x"60",x"00",x"37",x"00", -- 0x04A8
		x"75",x"00",x"76",x"00",x"77",x"00",x"39",x"00", -- 0x04B0
		x"75",x"00",x"74",x"00",x"76",x"00",x"77",x"00", -- 0x04B8
		x"77",x"00",x"74",x"00",x"75",x"00",x"76",x"00", -- 0x04C0
		x"74",x"00",x"3A",x"00",x"3B",x"00",x"75",x"00", -- 0x04C8
		x"3C",x"00",x"3D",x"00",x"3E",x"00",x"74",x"00", -- 0x04D0
		x"3F",x"00",x"70",x"00",x"40",x"00",x"75",x"00", -- 0x04D8
		x"51",x"80",x"50",x"80",x"61",x"00",x"76",x"00", -- 0x04E0
		x"53",x"80",x"2D",x"02",x"52",x"80",x"47",x"00", -- 0x04E8
		x"51",x"C0",x"44",x"C0",x"54",x"80",x"4B",x"00", -- 0x04F0
		x"71",x"00",x"56",x"80",x"54",x"C0",x"4B",x"00", -- 0x04F8
		x"72",x"00",x"59",x"40",x"52",x"C0",x"4A",x"00", -- 0x0500
		x"73",x"00",x"55",x"C0",x"33",x"00",x"74",x"00", -- 0x0508
		x"70",x"00",x"71",x"00",x"34",x"00",x"75",x"00", -- 0x0510
		x"5A",x"00",x"37",x"00",x"35",x"00",x"76",x"00", -- 0x0518
		x"75",x"00",x"39",x"00",x"77",x"00",x"74",x"00", -- 0x0520
		x"77",x"00",x"74",x"00",x"76",x"00",x"75",x"00", -- 0x0528
		x"75",x"00",x"76",x"00",x"75",x"00",x"76",x"00", -- 0x0530
		x"75",x"00",x"74",x"00",x"76",x"00",x"77",x"00", -- 0x0538
		x"77",x"00",x"74",x"00",x"75",x"00",x"76",x"00", -- 0x0540
		x"74",x"00",x"77",x"00",x"74",x"00",x"76",x"00", -- 0x0548
		x"77",x"00",x"76",x"00",x"77",x"00",x"75",x"00", -- 0x0550
		x"75",x"00",x"74",x"00",x"3C",x"00",x"3F",x"00", -- 0x0558
		x"77",x"00",x"3C",x"00",x"3F",x"00",x"55",x"00", -- 0x0560
		x"74",x"00",x"62",x"00",x"57",x"00",x"2D",x"02", -- 0x0568
		x"77",x"00",x"63",x"00",x"53",x"80",x"2D",x"02", -- 0x0570
		x"75",x"00",x"64",x"00",x"58",x"00",x"2D",x"02", -- 0x0578
		x"75",x"00",x"64",x"00",x"59",x"00",x"2D",x"02", -- 0x0580
		x"76",x"00",x"65",x"00",x"59",x"40",x"2D",x"02", -- 0x0588
		x"77",x"00",x"5C",x"00",x"5D",x"00",x"5D",x"80", -- 0x0590
		x"75",x"00",x"5E",x"00",x"5F",x"00",x"5F",x"80", -- 0x0598
		x"77",x"00",x"74",x"00",x"60",x"00",x"37",x"00", -- 0x05A0
		x"74",x"00",x"75",x"00",x"76",x"00",x"39",x"00", -- 0x05A8
		x"77",x"00",x"76",x"00",x"75",x"00",x"74",x"00", -- 0x05B0
		x"FF",x"FF",x"75",x"00",x"74",x"00",x"76",x"00", -- 0x05B8
		x"77",x"00",x"77",x"00",x"3A",x"00",x"3B",x"00", -- 0x05C0
		x"76",x"00",x"74",x"00",x"63",x"00",x"69",x"00", -- 0x05C8
		x"75",x"00",x"76",x"00",x"64",x"00",x"6A",x"00", -- 0x05D0
		x"74",x"00",x"75",x"00",x"68",x"00",x"6B",x"00", -- 0x05D8
		x"3F",x"00",x"66",x"00",x"67",x"00",x"31",x"40", -- 0x05E0
		x"32",x"40",x"70",x"00",x"71",x"00",x"2F",x"40", -- 0x05E8
		x"2A",x"40",x"2E",x"40",x"32",x"C0",x"2A",x"C0", -- 0x05F0
		x"6E",x"00",x"2A",x"40",x"2A",x"C0",x"6F",x"00", -- 0x05F8
		x"6D",x"00",x"6D",x"00",x"33",x"02",x"2C",x"00", -- 0x0600
		x"6E",x"00",x"6D",x"00",x"27",x"40",x"29",x"C0", -- 0x0608
		x"6F",x"00",x"24",x"40",x"00",x"00",x"27",x"C0", -- 0x0610
		x"2C",x"C0",x"00",x"00",x"01",x"00",x"02",x"00", -- 0x0618
		x"24",x"40",x"01",x"00",x"03",x"00",x"02",x"00", -- 0x0620
		x"00",x"00",x"03",x"00",x"00",x"00",x"01",x"00", -- 0x0628
		x"02",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x0630
		x"01",x"00",x"FF",x"FF",x"01",x"00",x"02",x"00", -- 0x0638
		x"03",x"00",x"00",x"00",x"00",x"00",x"03",x"00", -- 0x0640
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0648
		x"00",x"00",x"03",x"00",x"24",x"00",x"01",x"00", -- 0x0650
		x"03",x"00",x"00",x"00",x"6D",x"00",x"27",x"00", -- 0x0658
		x"01",x"00",x"24",x"00",x"6E",x"00",x"38",x"02", -- 0x0660
		x"27",x"80",x"2C",x"80",x"6F",x"00",x"2C",x"00", -- 0x0668
		x"33",x"C2",x"6F",x"00",x"6E",x"00",x"6E",x"00", -- 0x0670
		x"71",x"00",x"70",x"00",x"6D",x"00",x"70",x"00", -- 0x0678
		x"72",x"00",x"71",x"00",x"71",x"00",x"70",x"00", -- 0x0680
		x"72",x"00",x"73",x"00",x"70",x"00",x"71",x"00", -- 0x0688
		x"73",x"00",x"2B",x"00",x"72",x"00",x"70",x"00", -- 0x0690
		x"33",x"00",x"75",x"00",x"73",x"00",x"71",x"00", -- 0x0698
		x"34",x"00",x"76",x"00",x"36",x"00",x"37",x"00", -- 0x06A0
		x"35",x"00",x"77",x"00",x"38",x"00",x"39",x"00", -- 0x06A8
		x"76",x"00",x"74",x"00",x"75",x"00",x"74",x"00", -- 0x06B0
		x"77",x"00",x"75",x"00",x"FF",x"FF",x"76",x"00", -- 0x06B8
		x"77",x"00",x"74",x"00",x"75",x"00",x"74",x"00", -- 0x06C0
		x"76",x"00",x"78",x"00",x"79",x"00",x"75",x"00", -- 0x06C8
		x"74",x"00",x"7A",x"00",x"7B",x"00",x"77",x"00", -- 0x06D0
		x"7C",x"00",x"7D",x"00",x"7E",x"00",x"76",x"00", -- 0x06D8
		x"7F",x"00",x"80",x"00",x"75",x"00",x"78",x"00", -- 0x06E0
		x"79",x"00",x"7E",x"00",x"77",x"00",x"81",x"00", -- 0x06E8
		x"82",x"00",x"77",x"00",x"76",x"00",x"80",x"00", -- 0x06F0
		x"75",x"00",x"76",x"00",x"74",x"00",x"76",x"00", -- 0x06F8
		x"77",x"00",x"74",x"00",x"75",x"00",x"74",x"00", -- 0x0700
		x"83",x"00",x"75",x"00",x"77",x"00",x"75",x"00", -- 0x0708
		x"84",x"00",x"85",x"00",x"76",x"00",x"77",x"00", -- 0x0710
		x"86",x"00",x"87",x"00",x"74",x"00",x"76",x"00", -- 0x0718
		x"88",x"00",x"89",x"00",x"8A",x"00",x"74",x"00", -- 0x0720
		x"76",x"00",x"8B",x"00",x"89",x"00",x"75",x"00", -- 0x0728
		x"74",x"00",x"77",x"00",x"8B",x"00",x"77",x"00", -- 0x0730
		x"75",x"00",x"76",x"00",x"74",x"00",x"76",x"00", -- 0x0738
		x"77",x"00",x"74",x"00",x"75",x"00",x"74",x"00", -- 0x0740
		x"3A",x"00",x"3B",x"00",x"77",x"00",x"3C",x"00", -- 0x0748
		x"3D",x"00",x"3E",x"00",x"76",x"00",x"3F",x"00", -- 0x0750
		x"8C",x"00",x"40",x"00",x"74",x"00",x"8D",x"00", -- 0x0758
		x"8E",x"00",x"8F",x"00",x"75",x"00",x"98",x"C0", -- 0x0760
		x"2E",x"02",x"90",x"00",x"47",x"00",x"2E",x"02", -- 0x0768
		x"2F",x"02",x"91",x"00",x"4B",x"00",x"2F",x"02", -- 0x0770
		x"2E",x"02",x"92",x"00",x"96",x"00",x"2E",x"02", -- 0x0778
		x"2F",x"02",x"93",x"00",x"66",x"00",x"2F",x"02", -- 0x0780
		x"2E",x"02",x"94",x"00",x"95",x"00",x"2E",x"02", -- 0x0788
		x"2F",x"02",x"2E",x"02",x"97",x"00",x"2F",x"02", -- 0x0790
		x"2E",x"02",x"94",x"40",x"95",x"40",x"2E",x"02", -- 0x0798
		x"2F",x"02",x"93",x"40",x"70",x"00",x"2F",x"02", -- 0x07A0
		x"2E",x"02",x"92",x"40",x"71",x"00",x"2E",x"02", -- 0x07A8
		x"2F",x"02",x"91",x"40",x"72",x"00",x"2F",x"02", -- 0x07B0
		x"98",x"00",x"8D",x"C0",x"2B",x"00",x"2E",x"02", -- 0x07B8
		x"99",x"00",x"33",x"00",x"75",x"00",x"2F",x"02", -- 0x07C0
		x"9A",x"00",x"A4",x"00",x"77",x"00",x"2E",x"02", -- 0x07C8
		x"9B",x"00",x"A1",x"00",x"76",x"00",x"2F",x"02", -- 0x07D0
		x"9C",x"00",x"A2",x"00",x"74",x"00",x"2E",x"02", -- 0x07D8
		x"92",x"00",x"A3",x"00",x"75",x"00",x"2F",x"02", -- 0x07E0
		x"9D",x"00",x"70",x"00",x"47",x"00",x"2E",x"02", -- 0x07E8
		x"92",x"40",x"71",x"00",x"4B",x"00",x"2F",x"02", -- 0x07F0
		x"9E",x"00",x"72",x"00",x"4A",x"00",x"A0",x"00", -- 0x07F8
		x"9F",x"00",x"33",x"00",x"75",x"00",x"70",x"00", -- 0x0800
		x"71",x"00",x"34",x"00",x"77",x"00",x"36",x"00", -- 0x0808
		x"37",x"00",x"35",x"00",x"76",x"00",x"38",x"00", -- 0x0810
		x"39",x"00",x"76",x"00",x"74",x"00",x"76",x"00", -- 0x0818
		x"77",x"00",x"74",x"00",x"75",x"00",x"74",x"00", -- 0x0820
		x"76",x"00",x"75",x"00",x"77",x"00",x"75",x"00", -- 0x0828
		x"74",x"00",x"77",x"00",x"76",x"00",x"77",x"00", -- 0x0830
		x"75",x"00",x"76",x"00",x"74",x"00",x"76",x"00", -- 0x0838
		x"77",x"00",x"74",x"00",x"75",x"00",x"74",x"00", -- 0x0840
		x"76",x"00",x"78",x"00",x"79",x"00",x"75",x"00", -- 0x0848
		x"74",x"00",x"7A",x"00",x"7B",x"00",x"77",x"00", -- 0x0850
		x"A5",x"00",x"7D",x"00",x"7E",x"00",x"76",x"00", -- 0x0858
		x"A6",x"00",x"A8",x"00",x"75",x"00",x"78",x"00", -- 0x0860
		x"A7",x"00",x"A9",x"00",x"77",x"00",x"81",x"00", -- 0x0868
		x"AA",x"00",x"AB",x"00",x"76",x"00",x"80",x"00", -- 0x0870
		x"75",x"00",x"AC",x"00",x"8A",x"00",x"76",x"00", -- 0x0878
		x"77",x"00",x"8B",x"00",x"89",x"00",x"74",x"00", -- 0x0880
		x"76",x"00",x"75",x"00",x"8B",x"00",x"75",x"00", -- 0x0888
		x"74",x"00",x"77",x"00",x"76",x"00",x"77",x"00", -- 0x0890
		x"75",x"00",x"76",x"00",x"74",x"00",x"76",x"00", -- 0x0898
		x"77",x"00",x"74",x"00",x"75",x"00",x"74",x"00", -- 0x08A0
		x"76",x"00",x"75",x"00",x"77",x"00",x"75",x"00", -- 0x08A8
		x"74",x"00",x"77",x"00",x"76",x"00",x"77",x"00", -- 0x08B0
		x"75",x"00",x"76",x"00",x"74",x"00",x"FF",x"FF", -- 0x08B8
		x"76",x"00",x"3A",x"00",x"3B",x"00",x"75",x"00", -- 0x08C0
		x"74",x"00",x"63",x"00",x"69",x"00",x"77",x"00", -- 0x08C8
		x"75",x"00",x"64",x"00",x"6A",x"00",x"76",x"00", -- 0x08D0
		x"77",x"00",x"68",x"00",x"6B",x"00",x"3F",x"00", -- 0x08D8
		x"66",x"00",x"67",x"00",x"71",x"00",x"72",x"00", -- 0x08E0
		x"70",x"00",x"72",x"00",x"70",x"00",x"73",x"00", -- 0x08E8
		x"71",x"00",x"70",x"00",x"72",x"00",x"71",x"00", -- 0x08F0
		x"2D",x"C0",x"6D",x"00",x"70",x"00",x"72",x"00", -- 0x08F8
		x"00",x"00",x"29",x"C0",x"6E",x"00",x"28",x"C0", -- 0x0900
		x"01",x"00",x"27",x"C0",x"2C",x"80",x"25",x"C0", -- 0x0908
		x"02",x"00",x"01",x"00",x"24",x"40",x"00",x"00", -- 0x0910
		x"03",x"00",x"00",x"00",x"02",x"00",x"01",x"00", -- 0x0918
		x"00",x"00",x"03",x"00",x"01",x"00",x"02",x"00", -- 0x0920
		x"01",x"00",x"02",x"00",x"00",x"00",x"03",x"00", -- 0x0928
		x"02",x"00",x"01",x"00",x"03",x"00",x"00",x"00", -- 0x0930
		x"03",x"00",x"00",x"00",x"02",x"00",x"01",x"00", -- 0x0938
		x"FF",x"FF",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x0940
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x0948
		x"03",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x0950
		x"00",x"00",x"18",x"00",x"19",x"00",x"AD",x"00", -- 0x0958
		x"01",x"00",x"1A",x"00",x"20",x"00",x"AE",x"00", -- 0x0960
		x"02",x"00",x"1B",x"00",x"21",x"00",x"AF",x"00", -- 0x0968
		x"03",x"00",x"1C",x"00",x"22",x"00",x"B0",x"00", -- 0x0970
		x"00",x"00",x"1D",x"00",x"1E",x"00",x"B1",x"00", -- 0x0978
		x"01",x"00",x"00",x"00",x"03",x"00",x"11",x"00", -- 0x0980
		x"02",x"00",x"01",x"00",x"14",x"00",x"00",x"00", -- 0x0988
		x"03",x"00",x"02",x"00",x"0E",x"00",x"03",x"00", -- 0x0990
		x"00",x"00",x"03",x"00",x"17",x"00",x"02",x"00", -- 0x0998
		x"01",x"00",x"00",x"00",x"B2",x"00",x"01",x"00", -- 0x09A0
		x"02",x"00",x"B3",x"00",x"B4",x"00",x"00",x"00", -- 0x09A8
		x"03",x"00",x"B5",x"00",x"B7",x"00",x"04",x"00", -- 0x09B0
		x"05",x"00",x"B6",x"00",x"B8",x"00",x"06",x"00", -- 0x09B8
		x"07",x"00",x"B9",x"00",x"BE",x"00",x"08",x"00", -- 0x09C0
		x"09",x"00",x"BA",x"00",x"22",x"00",x"0A",x"00", -- 0x09C8
		x"0B",x"00",x"BB",x"00",x"21",x"00",x"0C",x"00", -- 0x09D0
		x"0D",x"00",x"BC",x"00",x"BD",x"00",x"72",x"02", -- 0x09D8
		x"10",x"00",x"00",x"00",x"03",x"00",x"12",x"00", -- 0x09E0
		x"13",x"00",x"01",x"00",x"02",x"00",x"15",x"00", -- 0x09E8
		x"16",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x09F0
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x09F8
		x"01",x"00",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x0A00
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x0A08
		x"03",x"00",x"17",x"00",x"01",x"00",x"03",x"00", -- 0x0A10
		x"00",x"00",x"03",x"00",x"11",x"00",x"02",x"00", -- 0x0A18
		x"01",x"00",x"19",x"00",x"32",x"02",x"01",x"00", -- 0x0A20
		x"02",x"00",x"20",x"00",x"AF",x"00",x"00",x"00", -- 0x0A28
		x"03",x"00",x"22",x"00",x"B0",x"00",x"03",x"00", -- 0x0A30
		x"00",x"00",x"1E",x"00",x"B1",x"00",x"02",x"00", -- 0x0A38
		x"01",x"00",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x0A40
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x0A48
		x"03",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x0A50
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x0A58
		x"01",x"00",x"00",x"00",x"03",x"00",x"BF",x"00", -- 0x0A60
		x"C0",x"00",x"01",x"00",x"02",x"00",x"C1",x"00", -- 0x0A68
		x"CA",x"00",x"02",x"00",x"01",x"00",x"C2",x"00", -- 0x0A70
		x"CB",x"00",x"03",x"00",x"C3",x"00",x"CC",x"00", -- 0x0A78
		x"CD",x"00",x"00",x"00",x"C4",x"00",x"CE",x"00", -- 0x0A80
		x"CF",x"00",x"01",x"00",x"C5",x"00",x"D0",x"00", -- 0x0A88
		x"D1",x"00",x"02",x"00",x"C4",x"40",x"D2",x"00", -- 0x0A90
		x"D3",x"00",x"03",x"00",x"C3",x"40",x"D4",x"00", -- 0x0A98
		x"20",x"00",x"00",x"00",x"03",x"00",x"C6",x"00", -- 0x0AA0
		x"D5",x"00",x"01",x"00",x"02",x"00",x"C7",x"00", -- 0x0AA8
		x"D6",x"00",x"02",x"00",x"01",x"00",x"C8",x"00", -- 0x0AB0
		x"D7",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x0AB8
		x"C9",x"00",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x0AC0
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x0AC8
		x"03",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x0AD0
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x0AD8
		x"01",x"00",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x0AE0
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x0AE8
		x"03",x"00",x"02",x"00",x"01",x"00",x"14",x"00", -- 0x0AF0
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x0AF8
		x"01",x"00",x"00",x"00",x"03",x"00",x"17",x"00", -- 0x0B00
		x"02",x"00",x"01",x"00",x"BF",x"00",x"D8",x"00", -- 0x0B08
		x"D9",x"00",x"02",x"00",x"DA",x"00",x"DB",x"00", -- 0x0B10
		x"DC",x"00",x"03",x"00",x"DD",x"00",x"DE",x"00", -- 0x0B18
		x"E4",x"00",x"00",x"00",x"E0",x"00",x"13",x"00", -- 0x0B20
		x"02",x"00",x"01",x"00",x"DF",x"00",x"E2",x"00", -- 0x0B28
		x"03",x"00",x"02",x"00",x"E1",x"00",x"E3",x"00", -- 0x0B30
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x0B38
		x"01",x"00",x"FF",x"FF",x"00",x"00",x"03",x"00", -- 0x0B40
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x0B48
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x0B50
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x0B58
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x0B60
		x"01",x"00",x"24",x"00",x"01",x"00",x"02",x"00", -- 0x0B68
		x"A5",x"01",x"2C",x"80",x"02",x"00",x"01",x"00", -- 0x0B70
		x"A4",x"01",x"6D",x"00",x"24",x"00",x"00",x"00", -- 0x0B78
		x"A3",x"01",x"6E",x"00",x"2C",x"00",x"A1",x"01", -- 0x0B80
		x"A2",x"01",x"6D",x"00",x"6E",x"00",x"EB",x"00", -- 0x0B88
		x"2C",x"80",x"6E",x"00",x"6F",x"00",x"6D",x"00", -- 0x0B90
		x"6E",x"00",x"6F",x"00",x"6E",x"00",x"6F",x"00", -- 0x0B98
		x"6D",x"00",x"6E",x"00",x"6D",x"00",x"6E",x"00", -- 0x0BA0
		x"6F",x"00",x"6D",x"00",x"6E",x"00",x"6F",x"00", -- 0x0BA8
		x"6D",x"00",x"6E",x"00",x"6F",x"00",x"6D",x"00", -- 0x0BB0
		x"6E",x"00",x"6F",x"00",x"6E",x"00",x"6F",x"00", -- 0x0BB8
		x"6D",x"00",x"6E",x"00",x"FF",x"FF",x"6D",x"00", -- 0x0BC0
		x"6E",x"00",x"6F",x"00",x"6D",x"00",x"9B",x"01", -- 0x0BC8
		x"6F",x"00",x"9A",x"01",x"6E",x"00",x"6F",x"00", -- 0x0BD0
		x"6D",x"00",x"9B",x"01",x"6F",x"00",x"9F",x"01", -- 0x0BD8
		x"6F",x"00",x"6D",x"00",x"9E",x"01",x"9D",x"01", -- 0x0BE0
		x"6E",x"00",x"9A",x"01",x"6D",x"00",x"6E",x"00", -- 0x0BE8
		x"9A",x"01",x"9C",x"01",x"6E",x"00",x"9E",x"01", -- 0x0BF0
		x"6D",x"00",x"9D",x"01",x"6F",x"00",x"6E",x"00", -- 0x0BF8
		x"9B",x"01",x"9F",x"01",x"6E",x"00",x"6D",x"00", -- 0x0C00
		x"9D",x"01",x"9E",x"01",x"9E",x"01",x"6E",x"00", -- 0x0C08
		x"A0",x"01",x"9E",x"01",x"6E",x"00",x"6F",x"00", -- 0x0C10
		x"9C",x"01",x"9C",x"01",x"9B",x"01",x"6E",x"00", -- 0x0C18
		x"6F",x"00",x"6D",x"00",x"6E",x"00",x"6D",x"00", -- 0x0C20
		x"9A",x"01",x"6F",x"00",x"9E",x"01",x"6E",x"00", -- 0x0C28
		x"6F",x"00",x"9B",x"01",x"6E",x"00",x"6F",x"00", -- 0x0C30
		x"9C",x"01",x"6E",x"00",x"6F",x"00",x"6E",x"00", -- 0x0C38
		x"6F",x"00",x"6D",x"00",x"6E",x"00",x"6D",x"00", -- 0x0C40
		x"6E",x"00",x"9C",x"01",x"6D",x"00",x"6E",x"00", -- 0x0C48
		x"6F",x"00",x"9E",x"01",x"6E",x"00",x"2A",x"80", -- 0x0C50
		x"6D",x"00",x"6E",x"00",x"6F",x"00",x"32",x"80", -- 0x0C58
		x"2A",x"80",x"6D",x"00",x"9F",x"01",x"70",x"00", -- 0x0C60
		x"2F",x"00",x"6F",x"00",x"9E",x"01",x"71",x"00", -- 0x0C68
		x"31",x"00",x"2A",x"80",x"6E",x"00",x"09",x"01", -- 0x0C70
		x"AC",x"01",x"A6",x"01",x"6F",x"00",x"20",x"00", -- 0x0C78
		x"AD",x"01",x"A7",x"01",x"6E",x"00",x"21",x"00", -- 0x0C80
		x"EA",x"00",x"31",x"00",x"A8",x"01",x"22",x"00", -- 0x0C88
		x"0A",x"01",x"70",x"00",x"A9",x"01",x"23",x"00", -- 0x0C90
		x"AE",x"01",x"71",x"00",x"AA",x"01",x"20",x"00", -- 0x0C98
		x"0B",x"01",x"72",x"00",x"AB",x"01",x"21",x"00", -- 0x0CA0
		x"20",x"00",x"AF",x"01",x"70",x"00",x"22",x"00", -- 0x0CA8
		x"21",x"00",x"B0",x"01",x"71",x"00",x"23",x"00", -- 0x0CB0
		x"20",x"00",x"0A",x"01",x"72",x"00",x"20",x"00", -- 0x0CB8
		x"23",x"00",x"B1",x"01",x"73",x"00",x"21",x"00", -- 0x0CC0
		x"20",x"00",x"35",x"02",x"70",x"00",x"22",x"00", -- 0x0CC8
		x"21",x"00",x"B2",x"01",x"71",x"00",x"23",x"00", -- 0x0CD0
		x"20",x"00",x"B3",x"01",x"72",x"00",x"20",x"00", -- 0x0CD8
		x"0C",x"01",x"70",x"00",x"73",x"00",x"21",x"00", -- 0x0CE0
		x"B4",x"01",x"71",x"00",x"70",x"00",x"22",x"00", -- 0x0CE8
		x"35",x"02",x"72",x"00",x"71",x"00",x"23",x"00", -- 0x0CF0
		x"B5",x"01",x"B7",x"01",x"72",x"00",x"F1",x"00", -- 0x0CF8
		x"B6",x"01",x"9D",x"80",x"B8",x"01",x"70",x"00", -- 0x0D00
		x"71",x"00",x"92",x"C0",x"B9",x"01",x"71",x"00", -- 0x0D08
		x"73",x"00",x"BA",x"01",x"BB",x"01",x"72",x"00", -- 0x0D10
		x"BC",x"01",x"BD",x"01",x"B9",x"C1",x"73",x"00", -- 0x0D18
		x"BE",x"01",x"8E",x"80",x"BF",x"01",x"70",x"00", -- 0x0D20
		x"C0",x"01",x"2E",x"02",x"C1",x"01",x"71",x"00", -- 0x0D28
		x"95",x"C0",x"2F",x"02",x"97",x"00",x"72",x"00", -- 0x0D30
		x"70",x"00",x"C2",x"01",x"95",x"40",x"73",x"00", -- 0x0D38
		x"72",x"00",x"8C",x"40",x"70",x"00",x"70",x"00", -- 0x0D40
		x"71",x"00",x"72",x"00",x"73",x"00",x"BD",x"01", -- 0x0D48
		x"73",x"00",x"70",x"00",x"36",x"02",x"8E",x"80", -- 0x0D50
		x"C3",x"01",x"E8",x"00",x"20",x"00",x"2E",x"02", -- 0x0D58
		x"97",x"00",x"14",x"01",x"21",x"00",x"2F",x"02", -- 0x0D60
		x"95",x"40",x"C4",x"01",x"22",x"00",x"8C",x"40", -- 0x0D68
		x"73",x"00",x"C5",x"01",x"23",x"00",x"72",x"00", -- 0x0D70
		x"70",x"00",x"C6",x"01",x"20",x"00",x"73",x"00", -- 0x0D78
		x"72",x"00",x"C7",x"01",x"21",x"00",x"70",x"00", -- 0x0D80
		x"71",x"00",x"C8",x"01",x"22",x"00",x"71",x"00", -- 0x0D88
		x"73",x"00",x"C9",x"01",x"23",x"00",x"72",x"00", -- 0x0D90
		x"70",x"00",x"CA",x"01",x"CB",x"01",x"73",x"00", -- 0x0D98
		x"72",x"00",x"71",x"00",x"F1",x"00",x"71",x"00", -- 0x0DA0
		x"70",x"00",x"72",x"00",x"70",x"00",x"72",x"00", -- 0x0DA8
		x"32",x"C0",x"31",x"C0",x"71",x"00",x"30",x"C0", -- 0x0DB0
		x"2A",x"C0",x"2F",x"C0",x"2E",x"C0",x"6E",x"00", -- 0x0DB8
		x"6D",x"00",x"2A",x"40",x"2A",x"C0",x"FF",x"FF", -- 0x0DC0
		x"6D",x"00",x"6E",x"00",x"6F",x"00",x"6D",x"00", -- 0x0DC8
		x"6E",x"00",x"6F",x"00",x"6D",x"00",x"6E",x"00", -- 0x0DD0
		x"6F",x"00",x"6D",x"00",x"6E",x"00",x"6F",x"00", -- 0x0DD8
		x"6E",x"00",x"6F",x"00",x"6D",x"00",x"6E",x"00", -- 0x0DE0
		x"6D",x"00",x"6E",x"00",x"6F",x"00",x"6D",x"00", -- 0x0DE8
		x"6E",x"00",x"6F",x"00",x"6D",x"00",x"6E",x"00", -- 0x0DF0
		x"6F",x"00",x"6D",x"00",x"6E",x"00",x"6F",x"00", -- 0x0DF8
		x"6E",x"00",x"6F",x"00",x"6D",x"00",x"6E",x"00", -- 0x0E00
		x"6D",x"00",x"6E",x"00",x"6F",x"00",x"6D",x"00", -- 0x0E08
		x"2D",x"C0",x"6D",x"00",x"6D",x"00",x"6E",x"00", -- 0x0E10
		x"00",x"00",x"29",x"C0",x"6E",x"00",x"28",x"C0", -- 0x0E18
		x"01",x"00",x"27",x"C0",x"2C",x"80",x"25",x"C0", -- 0x0E20
		x"00",x"00",x"03",x"00",x"24",x"40",x"02",x"00", -- 0x0E28
		x"01",x"00",x"02",x"00",x"00",x"00",x"03",x"00", -- 0x0E30
		x"02",x"00",x"01",x"00",x"03",x"00",x"00",x"00", -- 0x0E38
		x"03",x"00",x"00",x"00",x"02",x"00",x"01",x"00", -- 0x0E40
		x"FF",x"FF",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x0E48
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x0E50
		x"03",x"00",x"02",x"00",x"01",x"00",x"03",x"00", -- 0x0E58
		x"00",x"00",x"03",x"00",x"00",x"00",x"02",x"00", -- 0x0E60
		x"01",x"00",x"00",x"00",x"03",x"00",x"01",x"00", -- 0x0E68
		x"02",x"00",x"01",x"00",x"02",x"00",x"00",x"00", -- 0x0E70
		x"03",x"00",x"B2",x"00",x"01",x"00",x"03",x"00", -- 0x0E78
		x"00",x"00",x"B4",x"00",x"00",x"00",x"02",x"00", -- 0x0E80
		x"01",x"00",x"B7",x"00",x"04",x"00",x"05",x"00", -- 0x0E88
		x"24",x"00",x"31",x"00",x"2A",x"80",x"EB",x"00", -- 0x0E90
		x"2C",x"80",x"71",x"00",x"2F",x"00",x"2A",x"00", -- 0x0E98
		x"30",x"00",x"72",x"00",x"31",x"00",x"32",x"00", -- 0x0EA0
		x"70",x"00",x"73",x"00",x"E5",x"00",x"71",x"00", -- 0x0EA8
		x"72",x"00",x"70",x"00",x"E6",x"00",x"E7",x"00", -- 0x0EB0
		x"73",x"00",x"E8",x"00",x"20",x"00",x"21",x"00", -- 0x0EB8
		x"E9",x"00",x"21",x"00",x"22",x"00",x"23",x"00", -- 0x0EC0
		x"EA",x"00",x"FF",x"FF",x"20",x"00",x"21",x"00", -- 0x0EC8
		x"22",x"00",x"23",x"00",x"21",x"00",x"23",x"00", -- 0x0ED0
		x"20",x"00",x"22",x"00",x"22",x"00",x"EC",x"00", -- 0x0ED8
		x"23",x"00",x"20",x"00",x"23",x"00",x"ED",x"00", -- 0x0EE0
		x"EE",x"00",x"18",x"01",x"EF",x"00",x"F0",x"00", -- 0x0EE8
		x"F1",x"00",x"F2",x"00",x"F3",x"00",x"72",x"00", -- 0x0EF0
		x"70",x"00",x"73",x"00",x"F4",x"00",x"71",x"00", -- 0x0EF8
		x"94",x"01",x"70",x"00",x"F5",x"00",x"F6",x"00", -- 0x0F00
		x"95",x"01",x"71",x"00",x"20",x"00",x"F7",x"00", -- 0x0F08
		x"71",x"00",x"96",x"01",x"21",x"00",x"F8",x"00", -- 0x0F10
		x"94",x"01",x"73",x"00",x"22",x"00",x"F9",x"00", -- 0x0F18
		x"97",x"01",x"95",x"01",x"23",x"00",x"FA",x"00", -- 0x0F20
		x"72",x"00",x"71",x"00",x"F1",x"00",x"F2",x"00", -- 0x0F28
		x"96",x"01",x"FB",x"00",x"71",x"00",x"72",x"00", -- 0x0F30
		x"32",x"C0",x"FC",x"00",x"72",x"00",x"98",x"01", -- 0x0F38
		x"FD",x"00",x"31",x"80",x"94",x"01",x"70",x"00", -- 0x0F40
		x"FE",x"00",x"71",x"00",x"70",x"00",x"04",x"81", -- 0x0F48
		x"04",x"41",x"72",x"00",x"71",x"00",x"00",x"01", -- 0x0F50
		x"70",x"00",x"95",x"01",x"72",x"00",x"01",x"01", -- 0x0F58
		x"73",x"00",x"95",x"01",x"2E",x"40",x"02",x"01", -- 0x0F60
		x"72",x"00",x"99",x"01",x"2A",x"40",x"03",x"01", -- 0x0F68
		x"04",x"01",x"96",x"01",x"0E",x"01",x"31",x"80", -- 0x0F70
		x"05",x"01",x"73",x"00",x"72",x"00",x"71",x"00", -- 0x0F78
		x"06",x"01",x"31",x"C0",x"73",x"00",x"98",x"01", -- 0x0F80
		x"32",x"80",x"07",x"01",x"70",x"00",x"96",x"01", -- 0x0F88
		x"71",x"00",x"08",x"01",x"94",x"01",x"72",x"00", -- 0x0F90
		x"95",x"01",x"73",x"00",x"09",x"01",x"F6",x"00", -- 0x0F98
		x"94",x"01",x"96",x"01",x"23",x"00",x"EA",x"00", -- 0x0FA0
		x"72",x"00",x"71",x"00",x"20",x"00",x"F5",x"00", -- 0x0FA8
		x"F6",x"00",x"72",x"00",x"21",x"00",x"22",x"00", -- 0x0FB0
		x"EA",x"00",x"95",x"01",x"22",x"00",x"21",x"00", -- 0x0FB8
		x"0A",x"01",x"70",x"00",x"23",x"00",x"20",x"00", -- 0x0FC0
		x"0B",x"01",x"71",x"00",x"20",x"00",x"23",x"00", -- 0x0FC8
		x"0C",x"01",x"72",x"00",x"21",x"00",x"22",x"00", -- 0x0FD0
		x"35",x"02",x"73",x"00",x"22",x"00",x"EF",x"00", -- 0x0FD8
		x"0D",x"01",x"70",x"00",x"23",x"00",x"F3",x"00", -- 0x0FE0
		x"72",x"00",x"71",x"00",x"20",x"00",x"F8",x"00", -- 0x0FE8
		x"71",x"00",x"72",x"00",x"22",x"00",x"F8",x"00", -- 0x0FF0
		x"70",x"00",x"73",x"00",x"21",x"00",x"F9",x"00", -- 0x0FF8
		x"98",x"01",x"70",x"00",x"23",x"00",x"FA",x"00", -- 0x1000
		x"72",x"00",x"71",x"00",x"F1",x"00",x"F2",x"00", -- 0x1008
		x"96",x"01",x"72",x"00",x"71",x"00",x"72",x"00", -- 0x1010
		x"70",x"00",x"95",x"01",x"72",x"00",x"71",x"00", -- 0x1018
		x"95",x"01",x"99",x"01",x"73",x"00",x"98",x"01", -- 0x1020
		x"94",x"01",x"96",x"01",x"70",x"00",x"96",x"01", -- 0x1028
		x"98",x"01",x"73",x"00",x"71",x"00",x"71",x"00", -- 0x1030
		x"96",x"01",x"73",x"00",x"72",x"00",x"94",x"01", -- 0x1038
		x"71",x"00",x"95",x"01",x"94",x"01",x"70",x"00", -- 0x1040
		x"72",x"00",x"32",x"C0",x"70",x"00",x"73",x"00", -- 0x1048
		x"71",x"00",x"FD",x"00",x"71",x"00",x"98",x"01", -- 0x1050
		x"70",x"00",x"FE",x"00",x"94",x"01",x"96",x"01", -- 0x1058
		x"04",x"81",x"04",x"41",x"73",x"00",x"70",x"00", -- 0x1060
		x"00",x"01",x"71",x"00",x"2E",x"40",x"32",x"C0", -- 0x1068
		x"0F",x"01",x"72",x"00",x"2A",x"40",x"30",x"02", -- 0x1070
		x"32",x"00",x"98",x"01",x"0E",x"01",x"32",x"00", -- 0x1078
		x"73",x"00",x"96",x"01",x"73",x"00",x"70",x"00", -- 0x1080
		x"98",x"01",x"94",x"01",x"70",x"00",x"94",x"01", -- 0x1088
		x"71",x"00",x"72",x"00",x"94",x"01",x"95",x"01", -- 0x1090
		x"10",x"01",x"F6",x"00",x"72",x"00",x"73",x"00", -- 0x1098
		x"11",x"01",x"EA",x"00",x"73",x"00",x"12",x"01", -- 0x10A0
		x"13",x"01",x"21",x"00",x"70",x"00",x"14",x"01", -- 0x10A8
		x"21",x"00",x"22",x"00",x"71",x"00",x"E6",x"00", -- 0x10B0
		x"20",x"00",x"23",x"00",x"E8",x"00",x"21",x"00", -- 0x10B8
		x"23",x"00",x"20",x"00",x"23",x"00",x"20",x"00", -- 0x10C0
		x"22",x"00",x"21",x"00",x"FF",x"FF",x"20",x"00", -- 0x10C8
		x"23",x"00",x"21",x"00",x"22",x"00",x"21",x"00", -- 0x10D0
		x"22",x"00",x"20",x"00",x"23",x"00",x"22",x"00", -- 0x10D8
		x"21",x"00",x"23",x"00",x"20",x"00",x"23",x"00", -- 0x10E0
		x"20",x"00",x"22",x"00",x"21",x"00",x"15",x"01", -- 0x10E8
		x"21",x"00",x"21",x"00",x"22",x"00",x"16",x"01", -- 0x10F0
		x"22",x"00",x"20",x"00",x"23",x"00",x"BC",x"00", -- 0x10F8
		x"BD",x"00",x"0F",x"00",x"20",x"00",x"00",x"00", -- 0x1100
		x"01",x"00",x"12",x"00",x"21",x"00",x"00",x"00", -- 0x1108
		x"03",x"00",x"15",x"00",x"17",x"01",x"01",x"00", -- 0x1110
		x"02",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1118
		x"01",x"00",x"03",x"00",x"00",x"00",x"01",x"00", -- 0x1120
		x"00",x"00",x"02",x"00",x"01",x"00",x"00",x"00", -- 0x1128
		x"03",x"00",x"01",x"00",x"02",x"00",x"01",x"00", -- 0x1130
		x"02",x"00",x"00",x"00",x"03",x"00",x"02",x"00", -- 0x1138
		x"01",x"00",x"03",x"00",x"00",x"00",x"03",x"00", -- 0x1140
		x"00",x"00",x"02",x"00",x"01",x"00",x"FF",x"FF", -- 0x1148
		x"00",x"00",x"03",x"00",x"01",x"00",x"02",x"00", -- 0x1150
		x"01",x"00",x"02",x"00",x"00",x"00",x"03",x"00", -- 0x1158
		x"02",x"00",x"01",x"00",x"03",x"00",x"00",x"00", -- 0x1160
		x"03",x"00",x"00",x"00",x"02",x"00",x"01",x"00", -- 0x1168
		x"24",x"80",x"03",x"00",x"01",x"00",x"02",x"00", -- 0x1170
		x"2C",x"00",x"A5",x"81",x"00",x"00",x"03",x"00", -- 0x1178
		x"6D",x"00",x"A4",x"81",x"03",x"00",x"00",x"00", -- 0x1180
		x"6E",x"00",x"A3",x"81",x"02",x"00",x"24",x"80", -- 0x1188
		x"6F",x"00",x"A2",x"81",x"A1",x"81",x"2C",x"80", -- 0x1190
		x"6D",x"00",x"2C",x"00",x"EB",x"80",x"2A",x"00", -- 0x1198
		x"2A",x"00",x"2A",x"80",x"2A",x"00",x"32",x"00", -- 0x11A0
		x"32",x"00",x"32",x"80",x"32",x"00",x"70",x"00", -- 0x11A8
		x"70",x"00",x"CC",x"01",x"71",x"00",x"72",x"00", -- 0x11B0
		x"E8",x"00",x"CD",x"01",x"70",x"00",x"73",x"00", -- 0x11B8
		x"22",x"00",x"21",x"00",x"E7",x"00",x"70",x"00", -- 0x11C0
		x"23",x"00",x"20",x"00",x"22",x"00",x"E7",x"00", -- 0x11C8
		x"FF",x"FF",x"20",x"00",x"23",x"00",x"21",x"00", -- 0x11D0
		x"22",x"00",x"21",x"00",x"22",x"00",x"20",x"00", -- 0x11D8
		x"23",x"00",x"22",x"00",x"EC",x"00",x"23",x"00", -- 0x11E0
		x"20",x"00",x"F1",x"00",x"F2",x"00",x"EE",x"00", -- 0x11E8
		x"21",x"00",x"70",x"00",x"73",x"00",x"CE",x"01", -- 0x11F0
		x"22",x"00",x"71",x"00",x"72",x"00",x"37",x"02", -- 0x11F8
		x"23",x"00",x"B7",x"01",x"71",x"00",x"CF",x"01", -- 0x1200
		x"0D",x"01",x"D0",x"01",x"D1",x"01",x"72",x"00", -- 0x1208
		x"71",x"00",x"70",x"00",x"D2",x"01",x"71",x"00", -- 0x1210
		x"72",x"00",x"71",x"00",x"D3",x"01",x"D4",x"01", -- 0x1218
		x"73",x"00",x"F8",x"01",x"D5",x"01",x"D6",x"01", -- 0x1220
		x"70",x"00",x"F9",x"01",x"FA",x"01",x"D7",x"01", -- 0x1228
		x"71",x"00",x"FB",x"01",x"FC",x"01",x"D8",x"01", -- 0x1230
		x"72",x"00",x"FD",x"01",x"D9",x"01",x"DA",x"01", -- 0x1238
		x"73",x"00",x"72",x"00",x"DB",x"01",x"D4",x"41", -- 0x1240
		x"70",x"00",x"73",x"00",x"D8",x"C1",x"FE",x"01", -- 0x1248
		x"00",x"02",x"70",x"00",x"DC",x"01",x"01",x"02", -- 0x1250
		x"02",x"02",x"71",x"00",x"DD",x"01",x"03",x"02", -- 0x1258
		x"04",x"02",x"72",x"00",x"DE",x"01",x"05",x"02", -- 0x1260
		x"06",x"02",x"73",x"00",x"DE",x"41",x"07",x"02", -- 0x1268
		x"08",x"02",x"70",x"00",x"DD",x"41",x"71",x"00", -- 0x1270
		x"09",x"02",x"71",x"00",x"DF",x"01",x"72",x"00", -- 0x1278
		x"73",x"00",x"72",x"00",x"D3",x"01",x"E0",x"01", -- 0x1280
		x"01",x"02",x"73",x"00",x"E1",x"01",x"E2",x"01", -- 0x1288
		x"03",x"02",x"0A",x"02",x"72",x"00",x"E3",x"01", -- 0x1290
		x"05",x"02",x"0B",x"02",x"0C",x"02",x"DC",x"81", -- 0x1298
		x"07",x"02",x"0D",x"02",x"0E",x"02",x"DD",x"81", -- 0x12A0
		x"70",x"00",x"0F",x"02",x"10",x"02",x"E4",x"01", -- 0x12A8
		x"71",x"00",x"11",x"02",x"12",x"02",x"E5",x"01", -- 0x12B0
		x"72",x"00",x"13",x"02",x"72",x"00",x"E6",x"01", -- 0x12B8
		x"00",x"02",x"72",x"00",x"E1",x"41",x"E7",x"01", -- 0x12C0
		x"02",x"02",x"0C",x"02",x"D3",x"41",x"E8",x"01", -- 0x12C8
		x"04",x"02",x"0E",x"02",x"E3",x"81",x"05",x"02", -- 0x12D0
		x"06",x"02",x"10",x"02",x"E9",x"01",x"07",x"02", -- 0x12D8
		x"08",x"02",x"12",x"02",x"E9",x"01",x"73",x"00", -- 0x12E0
		x"09",x"02",x"14",x"02",x"EA",x"01",x"D5",x"C1", -- 0x12E8
		x"71",x"00",x"15",x"02",x"EB",x"01",x"EC",x"01", -- 0x12F0
		x"EC",x"81",x"16",x"02",x"17",x"02",x"ED",x"01", -- 0x12F8
		x"EE",x"01",x"18",x"02",x"19",x"02",x"EF",x"01", -- 0x1300
		x"8D",x"C0",x"1A",x"02",x"1B",x"02",x"F0",x"01", -- 0x1308
		x"72",x"00",x"1C",x"02",x"73",x"00",x"F1",x"01", -- 0x1310
		x"72",x"00",x"71",x"00",x"72",x"00",x"F2",x"01", -- 0x1318
		x"73",x"00",x"72",x"00",x"71",x"00",x"F3",x"01", -- 0x1320
		x"D5",x"C1",x"73",x"00",x"70",x"00",x"F4",x"01", -- 0x1328
		x"E2",x"01",x"70",x"00",x"73",x"00",x"71",x"00", -- 0x1330
		x"E3",x"01",x"1D",x"02",x"0A",x"02",x"70",x"00", -- 0x1338
		x"E9",x"81",x"1E",x"02",x"0B",x"02",x"0C",x"02", -- 0x1340
		x"F5",x"01",x"1F",x"02",x"0D",x"02",x"0E",x"02", -- 0x1348
		x"F6",x"01",x"20",x"02",x"0F",x"02",x"10",x"02", -- 0x1350
		x"72",x"00",x"21",x"02",x"11",x"02",x"12",x"02", -- 0x1358
		x"73",x"00",x"22",x"02",x"13",x"02",x"73",x"00", -- 0x1360
		x"70",x"00",x"73",x"00",x"70",x"00",x"72",x"00", -- 0x1368
		x"71",x"00",x"70",x"00",x"1D",x"02",x"0A",x"02", -- 0x1370
		x"72",x"00",x"23",x"02",x"1E",x"02",x"0B",x"02", -- 0x1378
		x"0C",x"02",x"24",x"02",x"1F",x"02",x"0D",x"02", -- 0x1380
		x"0E",x"02",x"25",x"02",x"20",x"02",x"0F",x"02", -- 0x1388
		x"10",x"02",x"26",x"02",x"21",x"02",x"11",x"02", -- 0x1390
		x"12",x"02",x"71",x"00",x"22",x"02",x"13",x"02", -- 0x1398
		x"73",x"00",x"72",x"00",x"71",x"00",x"73",x"00", -- 0x13A0
		x"70",x"00",x"09",x"01",x"AC",x"01",x"72",x"00", -- 0x13A8
		x"71",x"00",x"20",x"00",x"AD",x"01",x"71",x"00", -- 0x13B0
		x"72",x"00",x"21",x"00",x"F7",x"01",x"70",x"00", -- 0x13B8
		x"73",x"00",x"22",x"00",x"21",x"00",x"E7",x"00", -- 0x13C0
		x"70",x"00",x"23",x"00",x"20",x"00",x"22",x"00", -- 0x13C8
		x"E7",x"00",x"FF",x"FF",x"20",x"00",x"23",x"00", -- 0x13D0
		x"21",x"00",x"22",x"00",x"21",x"00",x"22",x"00", -- 0x13D8
		x"20",x"00",x"23",x"00",x"22",x"00",x"21",x"00", -- 0x13E0
		x"23",x"00",x"20",x"00",x"23",x"00",x"20",x"00", -- 0x13E8
		x"22",x"00",x"21",x"00",x"20",x"00",x"23",x"00", -- 0x13F0
		x"21",x"00",x"22",x"00",x"21",x"00",x"22",x"00", -- 0x13F8
		x"20",x"00",x"23",x"00",x"22",x"00",x"21",x"00", -- 0x1400
		x"23",x"00",x"20",x"00",x"12",x"00",x"20",x"00", -- 0x1408
		x"22",x"00",x"21",x"00",x"15",x"00",x"15",x"01", -- 0x1410
		x"21",x"00",x"22",x"00",x"01",x"00",x"16",x"01", -- 0x1418
		x"20",x"00",x"23",x"00",x"02",x"00",x"BC",x"00", -- 0x1420
		x"BD",x"00",x"17",x"01",x"03",x"00",x"00",x"00", -- 0x1428
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1430
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1438
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1440
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1448
		x"02",x"00",x"01",x"00",x"FF",x"FF",x"00",x"00", -- 0x1450
		x"03",x"00",x"01",x"00",x"02",x"00",x"7D",x"01", -- 0x1458
		x"7E",x"01",x"00",x"00",x"03",x"00",x"7F",x"01", -- 0x1460
		x"80",x"01",x"03",x"00",x"81",x"01",x"82",x"01", -- 0x1468
		x"83",x"01",x"84",x"01",x"83",x"01",x"85",x"01", -- 0x1470
		x"86",x"01",x"87",x"01",x"7F",x"01",x"88",x"01", -- 0x1478
		x"7F",x"01",x"83",x"01",x"86",x"01",x"82",x"01", -- 0x1480
		x"89",x"01",x"88",x"01",x"82",x"01",x"20",x"01", -- 0x1488
		x"1C",x"01",x"7F",x"01",x"1D",x"01",x"47",x"01", -- 0x1490
		x"23",x"01",x"24",x"01",x"25",x"01",x"26",x"01", -- 0x1498
		x"27",x"01",x"28",x"01",x"29",x"01",x"8B",x"01", -- 0x14A0
		x"2B",x"01",x"2C",x"01",x"35",x"01",x"8C",x"01", -- 0x14A8
		x"2F",x"01",x"8A",x"01",x"47",x"01",x"8D",x"01", -- 0x14B0
		x"8E",x"01",x"7A",x"01",x"1C",x"01",x"8F",x"01", -- 0x14B8
		x"90",x"01",x"66",x"01",x"91",x"01",x"72",x"00", -- 0x14C0
		x"92",x"01",x"6A",x"01",x"70",x"00",x"73",x"00", -- 0x14C8
		x"93",x"01",x"74",x"01",x"71",x"00",x"FF",x"FF", -- 0x14D0
		x"70",x"00",x"73",x"00",x"71",x"00",x"72",x"00", -- 0x14D8
		x"71",x"00",x"72",x"00",x"10",x"01",x"F6",x"00", -- 0x14E0
		x"72",x"00",x"70",x"00",x"11",x"01",x"27",x"02", -- 0x14E8
		x"73",x"00",x"12",x"01",x"13",x"01",x"21",x"00", -- 0x14F0
		x"70",x"00",x"14",x"01",x"21",x"00",x"22",x"00", -- 0x14F8
		x"71",x"00",x"E6",x"00",x"20",x"00",x"23",x"00", -- 0x1500
		x"72",x"00",x"28",x"02",x"23",x"00",x"18",x"01", -- 0x1508
		x"73",x"00",x"29",x"02",x"73",x"02",x"F2",x"00", -- 0x1510
		x"70",x"00",x"F1",x"00",x"F2",x"00",x"72",x"00", -- 0x1518
		x"71",x"00",x"72",x"00",x"70",x"00",x"73",x"00", -- 0x1520
		x"72",x"00",x"71",x"00",x"73",x"00",x"70",x"00", -- 0x1528
		x"73",x"00",x"76",x"01",x"72",x"00",x"71",x"00", -- 0x1530
		x"19",x"01",x"1A",x"01",x"71",x"00",x"74",x"01", -- 0x1538
		x"1B",x"01",x"1C",x"01",x"78",x"01",x"1D",x"01", -- 0x1540
		x"1E",x"01",x"1F",x"01",x"20",x"01",x"21",x"01", -- 0x1548
		x"22",x"01",x"23",x"01",x"24",x"01",x"25",x"01", -- 0x1550
		x"26",x"01",x"27",x"01",x"28",x"01",x"29",x"01", -- 0x1558
		x"2A",x"01",x"2B",x"01",x"2C",x"01",x"2D",x"01", -- 0x1560
		x"2E",x"01",x"2F",x"01",x"30",x"01",x"31",x"01", -- 0x1568
		x"32",x"01",x"33",x"01",x"34",x"01",x"35",x"01", -- 0x1570
		x"36",x"01",x"37",x"01",x"38",x"01",x"39",x"01", -- 0x1578
		x"2D",x"01",x"3B",x"01",x"3C",x"01",x"3D",x"01", -- 0x1580
		x"3E",x"01",x"3F",x"01",x"40",x"01",x"41",x"01", -- 0x1588
		x"42",x"01",x"43",x"01",x"44",x"01",x"45",x"01", -- 0x1590
		x"46",x"01",x"47",x"01",x"48",x"01",x"49",x"01", -- 0x1598
		x"4A",x"01",x"4B",x"01",x"4C",x"01",x"4D",x"01", -- 0x15A0
		x"4E",x"01",x"4F",x"01",x"50",x"01",x"51",x"01", -- 0x15A8
		x"52",x"01",x"53",x"01",x"54",x"01",x"55",x"01", -- 0x15B0
		x"56",x"01",x"57",x"01",x"58",x"01",x"59",x"01", -- 0x15B8
		x"5A",x"01",x"5B",x"01",x"5C",x"01",x"5D",x"01", -- 0x15C0
		x"5E",x"01",x"5F",x"01",x"60",x"01",x"61",x"01", -- 0x15C8
		x"62",x"01",x"3A",x"01",x"63",x"01",x"64",x"01", -- 0x15D0
		x"65",x"01",x"66",x"01",x"67",x"01",x"68",x"01", -- 0x15D8
		x"69",x"01",x"6A",x"01",x"6B",x"01",x"6C",x"01", -- 0x15E0
		x"6D",x"01",x"72",x"01",x"6E",x"01",x"6F",x"01", -- 0x15E8
		x"73",x"01",x"74",x"01",x"70",x"01",x"71",x"01", -- 0x15F0
		x"70",x"00",x"73",x"00",x"75",x"01",x"76",x"01", -- 0x15F8
		x"71",x"00",x"E5",x"00",x"77",x"01",x"78",x"01", -- 0x1600
		x"70",x"00",x"E6",x"00",x"E9",x"00",x"70",x"00", -- 0x1608
		x"E8",x"00",x"22",x"00",x"EA",x"00",x"71",x"00", -- 0x1610
		x"20",x"00",x"23",x"00",x"0A",x"01",x"72",x"00", -- 0x1618
		x"21",x"00",x"22",x"00",x"0B",x"01",x"73",x"00", -- 0x1620
		x"22",x"00",x"EC",x"00",x"0C",x"01",x"70",x"00", -- 0x1628
		x"23",x"00",x"ED",x"00",x"2A",x"02",x"71",x"00", -- 0x1630
		x"F1",x"00",x"F0",x"00",x"71",x"00",x"72",x"00", -- 0x1638
		x"71",x"00",x"72",x"00",x"70",x"00",x"73",x"00", -- 0x1640
		x"72",x"00",x"71",x"00",x"73",x"00",x"70",x"00", -- 0x1648
		x"73",x"00",x"70",x"00",x"72",x"00",x"71",x"00", -- 0x1650
		x"70",x"00",x"73",x"00",x"71",x"00",x"72",x"00", -- 0x1658
		x"71",x"00",x"1D",x"01",x"20",x"01",x"73",x"00", -- 0x1660
		x"19",x"01",x"79",x"01",x"7B",x"01",x"70",x"00", -- 0x1668
		x"1B",x"01",x"7A",x"01",x"1C",x"01",x"71",x"00", -- 0x1670
		x"1E",x"01",x"47",x"01",x"1F",x"01",x"1A",x"01", -- 0x1678
		x"22",x"01",x"23",x"01",x"47",x"01",x"52",x"01", -- 0x1680
		x"26",x"01",x"27",x"01",x"28",x"01",x"29",x"01", -- 0x1688
		x"2A",x"01",x"2B",x"01",x"2C",x"01",x"35",x"01", -- 0x1690
		x"2E",x"01",x"2F",x"01",x"7C",x"01",x"39",x"01", -- 0x1698
		x"32",x"01",x"3B",x"01",x"3C",x"01",x"3D",x"01", -- 0x16A0
		x"4F",x"01",x"3F",x"01",x"40",x"01",x"41",x"01", -- 0x16A8
		x"42",x"01",x"43",x"01",x"44",x"01",x"45",x"01", -- 0x16B0
		x"46",x"01",x"47",x"01",x"48",x"01",x"49",x"01", -- 0x16B8
		x"6D",x"01",x"6E",x"01",x"4C",x"01",x"4D",x"01", -- 0x16C0
		x"73",x"01",x"70",x"01",x"6E",x"01",x"1C",x"01", -- 0x16C8
		x"77",x"01",x"75",x"01",x"70",x"01",x"6A",x"01", -- 0x16D0
		x"FF",x"FF",x"70",x"00",x"73",x"00",x"77",x"01", -- 0x16D8
		x"78",x"01",x"71",x"00",x"72",x"00",x"70",x"00", -- 0x16E0
		x"73",x"00",x"72",x"00",x"71",x"00",x"73",x"00", -- 0x16E8
		x"70",x"00",x"E7",x"00",x"70",x"00",x"10",x"01", -- 0x16F0
		x"F6",x"00",x"20",x"00",x"E9",x"00",x"11",x"01", -- 0x16F8
		x"EA",x"00",x"21",x"00",x"F7",x"00",x"14",x"01", -- 0x1700
		x"23",x"00",x"22",x"00",x"F8",x"00",x"31",x"02", -- 0x1708
		x"20",x"00",x"23",x"00",x"F9",x"00",x"29",x"02", -- 0x1710
		x"21",x"00",x"20",x"00",x"FA",x"00",x"F1",x"00", -- 0x1718
		x"2B",x"02",x"F1",x"00",x"F2",x"00",x"70",x"00", -- 0x1720
		x"F1",x"00",x"72",x"00",x"32",x"C0",x"31",x"C0", -- 0x1728
		x"71",x"00",x"30",x"C0",x"2A",x"C0",x"2F",x"C0", -- 0x1730
		x"2E",x"C0",x"2D",x"C0",x"6D",x"00",x"2A",x"40", -- 0x1738
		x"2A",x"C0",x"01",x"00",x"29",x"C0",x"6E",x"00", -- 0x1740
		x"28",x"C0",x"02",x"00",x"27",x"C0",x"2C",x"80", -- 0x1748
		x"25",x"C0",x"03",x"00",x"00",x"00",x"24",x"40", -- 0x1750
		x"01",x"00",x"FF",x"FF",x"00",x"00",x"03",x"00", -- 0x1758
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1760
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1768
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1770
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1778
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1780
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1788
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1790
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1798
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x17A0
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x17A8
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x17B0
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x17B8
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x17C0
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x17C8
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x17D0
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x17D8
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x17E0
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x17E8
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x17F0
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x17F8
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1800
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1808
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1810
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1818
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1820
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1828
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1830
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1838
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1840
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1848
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1850
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1858
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1860
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1868
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1870
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1878
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1880
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1888
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1890
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1898
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x18A0
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x18A8
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x18B0
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x18B8
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x18C0
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x18C8
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x18D0
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x18D8
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x18E0
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x18E8
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x18F0
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x18F8
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1900
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1908
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1910
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1918
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1920
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1928
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1930
		x"02",x"00",x"01",x"00",x"00",x"00",x"03",x"00", -- 0x1938
		x"01",x"00",x"02",x"00",x"01",x"00",x"02",x"00", -- 0x1940
		x"00",x"00",x"03",x"00",x"02",x"00",x"01",x"00", -- 0x1948
		x"03",x"00",x"00",x"00",x"03",x"00",x"00",x"00", -- 0x1950
		x"02",x"00",x"01",x"00",x"FF",x"FF",x"3C",x"87", -- 0x1958
		x"3D",x"87",x"3E",x"87",x"3F",x"87",x"3D",x"87", -- 0x1960
		x"3C",x"87",x"3F",x"87",x"3E",x"87",x"3E",x"87", -- 0x1968
		x"3F",x"87",x"3C",x"87",x"3D",x"87",x"3F",x"87", -- 0x1970
		x"3E",x"87",x"3D",x"87",x"3C",x"87",x"32",x"E1", -- 0x1978
		x"2F",x"A1",x"35",x"A1",x"2D",x"A1",x"36",x"E1", -- 0x1980
		x"27",x"C1",x"3C",x"87",x"3D",x"87",x"39",x"02", -- 0x1988
		x"2C",x"62",x"3C",x"02",x"3D",x"02",x"3D",x"02", -- 0x1990
		x"23",x"C1",x"3D",x"87",x"3C",x"87",x"2F",x"0A", -- 0x1998
		x"30",x"0A",x"2E",x"62",x"39",x"02",x"2D",x"62", -- 0x19A0
		x"21",x"E1",x"3F",x"87",x"3E",x"87",x"17",x"02", -- 0x19A8
		x"18",x"02",x"16",x"02",x"31",x"0A",x"29",x"62", -- 0x19B0
		x"3C",x"02",x"25",x"C1",x"3C",x"87",x"23",x"02", -- 0x19B8
		x"22",x"02",x"13",x"02",x"2F",x"0A",x"2F",x"0A", -- 0x19C0
		x"2A",x"62",x"20",x"E1",x"27",x"C1",x"3E",x"87", -- 0x19C8
		x"1D",x"89",x"3C",x"87",x"3D",x"87",x"00",x"89", -- 0x19D0
		x"22",x"02",x"23",x"02",x"24",x"02",x"18",x"02", -- 0x19D8
		x"15",x"02",x"2B",x"62",x"23",x"C1",x"1E",x"89", -- 0x19E0
		x"3C",x"87",x"3F",x"87",x"3E",x"87",x"01",x"89", -- 0x19E8
		x"07",x"89",x"00",x"89",x"22",x"02",x"23",x"02", -- 0x19F0
		x"24",x"02",x"3A",x"88",x"26",x"E1",x"3C",x"87", -- 0x19F8
		x"3D",x"87",x"1F",x"89",x"3C",x"87",x"3D",x"87", -- 0x1A00
		x"3C",x"87",x"01",x"89",x"07",x"89",x"02",x"89", -- 0x1A08
		x"03",x"89",x"0D",x"89",x"3D",x"87",x"3F",x"87", -- 0x1A10
		x"3E",x"87",x"3D",x"87",x"1E",x"89",x"3C",x"87", -- 0x1A18
		x"3D",x"87",x"3E",x"87",x"11",x"89",x"12",x"89", -- 0x1A20
		x"13",x"89",x"14",x"89",x"1C",x"89",x"3D",x"87", -- 0x1A28
		x"11",x"89",x"1C",x"89",x"0E",x"E9",x"3F",x"87", -- 0x1A30
		x"10",x"89",x"22",x"02",x"23",x"02",x"3E",x"87", -- 0x1A38
		x"18",x"89",x"24",x"02",x"25",x"02",x"3F",x"87", -- 0x1A40
		x"01",x"89",x"07",x"89",x"02",x"89",x"09",x"89", -- 0x1A48
		x"08",x"89",x"05",x"89",x"06",x"89",x"00",x"00", -- 0x1A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"22",x"02", -- 0x1A58
		x"23",x"02",x"24",x"02",x"25",x"02",x"23",x"02", -- 0x1A60
		x"22",x"02",x"25",x"02",x"24",x"02",x"25",x"02", -- 0x1A68
		x"24",x"02",x"23",x"02",x"22",x"02",x"24",x"02", -- 0x1A70
		x"25",x"02",x"22",x"02",x"23",x"02",x"38",x"81", -- 0x1A78
		x"2E",x"A1",x"2E",x"A1",x"38",x"C1",x"38",x"A1", -- 0x1A80
		x"27",x"81",x"2E",x"A1",x"31",x"A1",x"3A",x"02", -- 0x1A88
		x"3B",x"02",x"3C",x"02",x"3A",x"02",x"31",x"E1", -- 0x1A90
		x"2E",x"A1",x"27",x"C1",x"3C",x"87",x"00",x"00", -- 0x1A98
		x"20",x"A1",x"3B",x"02",x"3C",x"02",x"3D",x"02", -- 0x1AA0
		x"3E",x"02",x"20",x"E1",x"38",x"C1",x"3C",x"02", -- 0x1AA8
		x"3B",x"02",x"2C",x"22",x"39",x"02",x"CA",x"02", -- 0x1AB0
		x"D6",x"02",x"CC",x"02",x"00",x"87",x"3B",x"02", -- 0x1AB8
		x"3C",x"02",x"3D",x"02",x"3A",x"42",x"31",x"E1", -- 0x1AC0
		x"2E",x"A1",x"31",x"A1",x"00",x"00",x"00",x"00", -- 0x1AC8
		x"2E",x"22",x"2F",x"0A",x"30",x"0A",x"31",x"0A", -- 0x1AD0
		x"32",x"0A",x"2A",x"62",x"3B",x"02",x"39",x"02", -- 0x1AD8
		x"39",x"02",x"2C",x"62",x"2C",x"62",x"2F",x"0A", -- 0x1AE0
		x"30",x"0A",x"31",x"0A",x"2E",x"62",x"39",x"02", -- 0x1AE8
		x"2E",x"22",x"30",x"0A",x"31",x"0A",x"32",x"0A", -- 0x1AF0
		x"31",x"0A",x"2F",x"0A",x"CD",x"02",x"2F",x"0A", -- 0x1AF8
		x"CA",x"02",x"CC",x"02",x"DB",x"02",x"CD",x"02", -- 0x1B00
		x"DB",x"02",x"DC",x"02",x"DD",x"02",x"30",x"0A", -- 0x1B08
		x"31",x"0A",x"CA",x"02",x"D6",x"02",x"C0",x"02", -- 0x1B10
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"32",x"0A", -- 0x1B18
		x"CD",x"02",x"DB",x"02",x"DC",x"02",x"DB",x"02", -- 0x1B20
		x"C2",x"02",x"D6",x"02",x"CC",x"02",x"DB",x"02", -- 0x1B28
		x"DC",x"02",x"C7",x"02",x"D7",x"02",x"D7",x"02", -- 0x1B30
		x"D1",x"02",x"DB",x"02",x"DC",x"02",x"DB",x"02", -- 0x1B38
		x"DC",x"02",x"DD",x"02",x"C7",x"02",x"D7",x"02", -- 0x1B40
		x"C5",x"02",x"2F",x"0A",x"30",x"0A",x"31",x"0A", -- 0x1B48
		x"32",x"0A",x"D2",x"02",x"DB",x"02",x"D7",x"02", -- 0x1B50
		x"D7",x"02",x"C5",x"02",x"31",x"0A",x"2F",x"0A", -- 0x1B58
		x"30",x"0A",x"31",x"0A",x"D0",x"02",x"00",x"00", -- 0x1B60
		x"F9",x"23",x"FA",x"23",x"F8",x"63",x"2F",x"0A", -- 0x1B68
		x"30",x"0A",x"F9",x"23",x"FA",x"23",x"F9",x"63", -- 0x1B70
		x"31",x"0A",x"32",x"0A",x"D3",x"02",x"FD",x"03", -- 0x1B78
		x"FD",x"03",x"FD",x"03",x"F5",x"63",x"FA",x"23", -- 0x1B80
		x"F6",x"23",x"FC",x"23",x"FD",x"03",x"FD",x"03", -- 0x1B88
		x"FB",x"63",x"2F",x"0A",x"30",x"0A",x"D0",x"02", -- 0x1B90
		x"DB",x"02",x"DC",x"02",x"DD",x"02",x"FD",x"03", -- 0x1B98
		x"FB",x"43",x"31",x"0A",x"32",x"0A",x"F7",x"43", -- 0x1BA0
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"CB",x"02", -- 0x1BA8
		x"DC",x"02",x"DD",x"02",x"DB",x"02",x"D4",x"02", -- 0x1BB0
		x"DD",x"02",x"DB",x"02",x"DC",x"02",x"FD",x"03", -- 0x1BB8
		x"F6",x"43",x"FA",x"03",x"F9",x"43",x"00",x"00", -- 0x1BC0
		x"F9",x"03",x"FA",x"03",x"FA",x"03",x"F9",x"43", -- 0x1BC8
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"DB",x"02", -- 0x1BD0
		x"DC",x"02",x"C8",x"02",x"2F",x"0A",x"F9",x"23", -- 0x1BD8
		x"FA",x"23",x"FA",x"23",x"FA",x"23",x"F8",x"63", -- 0x1BE0
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"30",x"0A", -- 0x1BE8
		x"2F",x"0A",x"F8",x"23",x"F6",x"23",x"F3",x"43", -- 0x1BF0
		x"30",x"0A",x"31",x"0A",x"32",x"0A",x"2F",x"0A", -- 0x1BF8
		x"30",x"0A",x"F4",x"23",x"FD",x"03",x"F9",x"23", -- 0x1C00
		x"FA",x"23",x"F9",x"63",x"31",x"0A",x"FD",x"03", -- 0x1C08
		x"FD",x"03",x"FD",x"03",x"F3",x"43",x"2F",x"0A", -- 0x1C10
		x"30",x"0A",x"31",x"0A",x"FB",x"23",x"30",x"0A", -- 0x1C18
		x"F9",x"23",x"FA",x"23",x"F5",x"23",x"FB",x"23", -- 0x1C20
		x"FD",x"03",x"FD",x"03",x"FD",x"03",x"00",x"00", -- 0x1C28
		x"C2",x"02",x"D6",x"02",x"D6",x"02",x"DB",x"02", -- 0x1C30
		x"C3",x"02",x"2F",x"0A",x"30",x"0A",x"DC",x"02", -- 0x1C38
		x"DD",x"02",x"C3",x"02",x"31",x"0A",x"32",x"0A", -- 0x1C40
		x"F7",x"03",x"FD",x"03",x"FD",x"03",x"DB",x"02", -- 0x1C48
		x"DC",x"02",x"DD",x"02",x"C2",x"02",x"C0",x"02", -- 0x1C50
		x"2F",x"0A",x"F9",x"03",x"FA",x"03",x"DB",x"02", -- 0x1C58
		x"C2",x"02",x"D6",x"02",x"D6",x"02",x"2F",x"0A", -- 0x1C60
		x"30",x"0A",x"31",x"0A",x"D3",x"02",x"DB",x"02", -- 0x1C68
		x"DC",x"02",x"C8",x"02",x"2F",x"0A",x"DB",x"02", -- 0x1C70
		x"C6",x"02",x"30",x"0A",x"31",x"0A",x"DC",x"02", -- 0x1C78
		x"D5",x"02",x"2F",x"0A",x"30",x"0A",x"DD",x"02", -- 0x1C80
		x"C1",x"02",x"31",x"0A",x"32",x"0A",x"2F",x"0A", -- 0x1C88
		x"CF",x"02",x"D7",x"02",x"D7",x"02",x"C5",x"02", -- 0x1C90
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"DB",x"02", -- 0x1C98
		x"C9",x"02",x"2F",x"0A",x"30",x"0A",x"2F",x"0A", -- 0x1CA0
		x"30",x"0A",x"D0",x"02",x"DB",x"02",x"30",x"0A", -- 0x1CA8
		x"31",x"0A",x"D3",x"02",x"DC",x"02",x"31",x"0A", -- 0x1CB0
		x"32",x"0A",x"2F",x"0A",x"CF",x"02",x"3C",x"02", -- 0x1CB8
		x"3D",x"02",x"20",x"C1",x"31",x"81",x"3B",x"02", -- 0x1CC0
		x"3C",x"02",x"3D",x"02",x"3E",x"02",x"3D",x"02", -- 0x1CC8
		x"3E",x"02",x"3B",x"02",x"3C",x"02",x"3C",x"02", -- 0x1CD0
		x"3D",x"02",x"3E",x"02",x"3B",x"02",x"2F",x"0A", -- 0x1CD8
		x"30",x"0A",x"31",x"0A",x"32",x"0A",x"31",x"0A", -- 0x1CE0
		x"32",x"0A",x"2F",x"0A",x"30",x"0A",x"30",x"0A", -- 0x1CE8
		x"2F",x"0A",x"32",x"0A",x"31",x"0A",x"32",x"0A", -- 0x1CF0
		x"31",x"0A",x"30",x"0A",x"2F",x"0A",x"DB",x"02", -- 0x1CF8
		x"DC",x"02",x"DD",x"02",x"23",x"02",x"DC",x"02", -- 0x1D00
		x"22",x"02",x"DB",x"02",x"DD",x"02",x"DD",x"02", -- 0x1D08
		x"DB",x"02",x"24",x"02",x"DC",x"02",x"25",x"02", -- 0x1D10
		x"DD",x"02",x"DC",x"02",x"DB",x"02",x"DB",x"02", -- 0x1D18
		x"DC",x"02",x"C7",x"05",x"D7",x"05",x"D7",x"05", -- 0x1D20
		x"D7",x"05",x"C5",x"05",x"CA",x"05",x"C7",x"05", -- 0x1D28
		x"C5",x"05",x"DA",x"25",x"D8",x"05",x"DA",x"45", -- 0x1D30
		x"CA",x"05",x"D6",x"05",x"00",x"00",x"DB",x"02", -- 0x1D38
		x"DC",x"02",x"DD",x"02",x"C6",x"05",x"DA",x"25", -- 0x1D40
		x"D9",x"05",x"CA",x"05",x"D6",x"05",x"CC",x"05", -- 0x1D48
		x"DB",x"02",x"DC",x"02",x"DD",x"02",x"DC",x"02", -- 0x1D50
		x"DD",x"02",x"DB",x"02",x"C9",x"05",x"DA",x"45", -- 0x1D58
		x"CD",x"05",x"DB",x"02",x"DC",x"02",x"00",x"00", -- 0x1D60
		x"C5",x"05",x"CA",x"05",x"D6",x"05",x"D6",x"05", -- 0x1D68
		x"D6",x"05",x"CC",x"05",x"DB",x"02",x"DB",x"02", -- 0x1D70
		x"DC",x"02",x"C7",x"05",x"D1",x"05",x"DD",x"02", -- 0x1D78
		x"C6",x"05",x"DA",x"25",x"DA",x"65",x"D1",x"05", -- 0x1D80
		x"DB",x"02",x"DC",x"02",x"DD",x"02",x"DC",x"02", -- 0x1D88
		x"C1",x"05",x"DA",x"05",x"D8",x"05",x"DA",x"65", -- 0x1D90
		x"D2",x"05",x"DB",x"02",x"DC",x"02",x"DD",x"02", -- 0x1D98
		x"DB",x"02",x"C2",x"05",x"D6",x"05",x"C0",x"05", -- 0x1DA0
		x"DA",x"05",x"CF",x"05",x"D7",x"05",x"D7",x"05", -- 0x1DA8
		x"D1",x"05",x"DB",x"02",x"00",x"00",x"DB",x"02", -- 0x1DB0
		x"C2",x"05",x"D6",x"05",x"D6",x"05",x"2F",x"0A", -- 0x1DB8
		x"41",x"23",x"42",x"23",x"41",x"63",x"2F",x"0A", -- 0x1DC0
		x"30",x"0A",x"41",x"23",x"42",x"23",x"40",x"23", -- 0x1DC8
		x"49",x"23",x"4A",x"03",x"49",x"63",x"40",x"63", -- 0x1DD0
		x"44",x"63",x"2F",x"0A",x"D3",x"02",x"4B",x"03", -- 0x1DD8
		x"46",x"63",x"30",x"0A",x"31",x"0A",x"4A",x"03", -- 0x1DE0
		x"49",x"63",x"48",x"63",x"32",x"0A",x"4B",x"03", -- 0x1DE8
		x"4A",x"03",x"49",x"63",x"43",x"63",x"4A",x"03", -- 0x1DF0
		x"4B",x"03",x"4A",x"03",x"46",x"63",x"4B",x"03", -- 0x1DF8
		x"4A",x"03",x"4B",x"03",x"49",x"63",x"43",x"63", -- 0x1E00
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"D3",x"02", -- 0x1E08
		x"DB",x"02",x"DC",x"02",x"DD",x"02",x"45",x"43", -- 0x1E10
		x"31",x"0A",x"32",x"0A",x"2F",x"0A",x"4A",x"03", -- 0x1E18
		x"49",x"43",x"40",x"43",x"42",x"03",x"4B",x"03", -- 0x1E20
		x"46",x"43",x"2F",x"0A",x"30",x"0A",x"4A",x"03", -- 0x1E28
		x"45",x"43",x"31",x"0A",x"32",x"0A",x"4B",x"03", -- 0x1E30
		x"47",x"63",x"44",x"63",x"2F",x"0A",x"4A",x"03", -- 0x1E38
		x"4B",x"03",x"46",x"63",x"30",x"0A",x"4B",x"03", -- 0x1E40
		x"4A",x"03",x"4B",x"03",x"45",x"43",x"49",x"43", -- 0x1E48
		x"40",x"43",x"41",x"43",x"31",x"0A",x"41",x"43", -- 0x1E50
		x"2F",x"0A",x"30",x"0A",x"32",x"0A",x"2F",x"0A", -- 0x1E58
		x"41",x"03",x"42",x"03",x"42",x"03",x"2F",x"0A", -- 0x1E60
		x"30",x"0A",x"D4",x"02",x"DB",x"02",x"31",x"0A", -- 0x1E68
		x"32",x"0A",x"D3",x"02",x"DC",x"02",x"30",x"0A", -- 0x1E70
		x"2F",x"0A",x"31",x"0A",x"D2",x"02",x"31",x"0A", -- 0x1E78
		x"32",x"0A",x"CE",x"02",x"DD",x"02",x"DB",x"02", -- 0x1E80
		x"DC",x"02",x"DD",x"02",x"C8",x"05",x"DD",x"02", -- 0x1E88
		x"DB",x"02",x"C8",x"05",x"DA",x"25",x"D7",x"05", -- 0x1E90
		x"C5",x"05",x"CA",x"05",x"C0",x"05",x"D8",x"05", -- 0x1E98
		x"CE",x"05",x"DB",x"02",x"DC",x"02",x"DA",x"05", -- 0x1EA0
		x"D4",x"05",x"DD",x"02",x"DB",x"02",x"D6",x"05", -- 0x1EA8
		x"CC",x"05",x"DB",x"02",x"DC",x"02",x"C4",x"05", -- 0x1EB0
		x"D3",x"05",x"DC",x"05",x"DD",x"02",x"C1",x"05", -- 0x1EB8
		x"DA",x"05",x"CF",x"05",x"D7",x"05",x"15",x"89", -- 0x1EC0
		x"3C",x"87",x"3D",x"87",x"3C",x"87",x"16",x"89", -- 0x1EC8
		x"15",x"89",x"3C",x"87",x"3D",x"87",x"22",x"02", -- 0x1ED0
		x"1A",x"89",x"3D",x"87",x"3C",x"87",x"23",x"02", -- 0x1ED8
		x"18",x"C9",x"3C",x"87",x"3D",x"87",x"07",x"89", -- 0x1EE0
		x"0A",x"89",x"3C",x"87",x"3D",x"87",x"27",x"81", -- 0x1EE8
		x"36",x"A1",x"2D",x"A1",x"26",x"C1",x"3C",x"87", -- 0x1EF0
		x"3D",x"87",x"3C",x"87",x"27",x"81",x"20",x"A1", -- 0x1EF8
		x"3B",x"02",x"3C",x"02",x"21",x"E1",x"3C",x"87", -- 0x1F00
		x"3D",x"87",x"3C",x"87",x"21",x"A1",x"3C",x"87", -- 0x1F08
		x"3D",x"87",x"25",x"81",x"2B",x"02",x"2C",x"22", -- 0x1F10
		x"39",x"02",x"2C",x"62",x"3A",x"02",x"0A",x"02", -- 0x1F18
		x"18",x"02",x"15",x"02",x"2E",x"62",x"3C",x"87", -- 0x1F20
		x"3D",x"87",x"23",x"81",x"38",x"02",x"3C",x"87", -- 0x1F28
		x"3D",x"87",x"26",x"A1",x"39",x"88",x"3C",x"87", -- 0x1F30
		x"3D",x"87",x"3C",x"87",x"18",x"89",x"3C",x"87", -- 0x1F38
		x"3D",x"87",x"3C",x"87",x"01",x"89",x"02",x"89", -- 0x1F40
		x"03",x"89",x"09",x"89",x"07",x"89",x"07",x"02", -- 0x1F48
		x"22",x"02",x"23",x"02",x"14",x"02",x"3C",x"87", -- 0x1F50
		x"3D",x"87",x"3C",x"87",x"38",x"81",x"36",x"A1", -- 0x1F58
		x"2D",x"A1",x"36",x"E1",x"00",x"00",x"3C",x"87", -- 0x1F60
		x"38",x"81",x"31",x"A1",x"3A",x"02",x"33",x"A1", -- 0x1F68
		x"3A",x"02",x"3C",x"02",x"3D",x"02",x"3C",x"87", -- 0x1F70
		x"3D",x"87",x"3C",x"87",x"25",x"81",x"3C",x"87", -- 0x1F78
		x"3D",x"87",x"3C",x"87",x"22",x"A1",x"3C",x"87", -- 0x1F80
		x"3D",x"87",x"3C",x"87",x"28",x"81",x"33",x"81", -- 0x1F88
		x"3A",x"21",x"2A",x"02",x"03",x"02",x"3D",x"87", -- 0x1F90
		x"33",x"81",x"3A",x"21",x"2C",x"02",x"3C",x"87", -- 0x1F98
		x"3D",x"87",x"38",x"A1",x"31",x"81",x"38",x"A1", -- 0x1FA0
		x"36",x"81",x"2D",x"81",x"00",x"00",x"3B",x"02", -- 0x1FA8
		x"71",x"04",x"72",x"04",x"00",x"00",x"6E",x"04", -- 0x1FB0
		x"6F",x"04",x"70",x"04",x"00",x"00",x"3A",x"02", -- 0x1FB8
		x"2C",x"22",x"39",x"02",x"6A",x"04",x"6B",x"04", -- 0x1FC0
		x"6C",x"04",x"6D",x"04",x"00",x"00",x"2B",x"22", -- 0x1FC8
		x"0A",x"02",x"18",x"02",x"66",x"04",x"67",x"04", -- 0x1FD0
		x"68",x"04",x"69",x"04",x"00",x"00",x"38",x"02", -- 0x1FD8
		x"1B",x"02",x"22",x"02",x"23",x"02",x"63",x"04", -- 0x1FE0
		x"64",x"04",x"65",x"04",x"00",x"00",x"2B",x"02", -- 0x1FE8
		x"00",x"02",x"23",x"02",x"24",x"02",x"60",x"04", -- 0x1FF0
		x"61",x"04",x"62",x"04",x"00",x"00",x"3A",x"21", -- 0x1FF8
		x"2A",x"02",x"02",x"02",x"25",x"02",x"05",x"02", -- 0x2000
		x"22",x"02",x"23",x"02",x"24",x"02",x"2E",x"02", -- 0x2008
		x"03",x"02",x"19",x"02",x"00",x"00",x"3A",x"22", -- 0x2010
		x"2C",x"02",x"39",x"22",x"00",x"00",x"2E",x"A1", -- 0x2018
		x"2E",x"A1",x"31",x"A1",x"31",x"E1",x"27",x"C1", -- 0x2020
		x"3C",x"87",x"3C",x"87",x"3D",x"87",x"3C",x"87", -- 0x2028
		x"3D",x"87",x"33",x"A1",x"2C",x"22",x"39",x"02", -- 0x2030
		x"2C",x"62",x"3C",x"02",x"3D",x"02",x"23",x"C1", -- 0x2038
		x"3D",x"87",x"3C",x"87",x"3D",x"87",x"3C",x"87", -- 0x2040
		x"25",x"81",x"2B",x"22",x"0A",x"02",x"18",x"02", -- 0x2048
		x"15",x"02",x"2B",x"62",x"20",x"C1",x"3C",x"87", -- 0x2050
		x"26",x"A1",x"39",x"88",x"23",x"02",x"3C",x"87", -- 0x2058
		x"23",x"81",x"38",x"02",x"07",x"02",x"3D",x"87", -- 0x2060
		x"3D",x"87",x"0C",x"89",x"07",x"89",x"22",x"02", -- 0x2068
		x"0E",x"89",x"0A",x"89",x"3D",x"87",x"07",x"89", -- 0x2070
		x"0A",x"89",x"3C",x"87",x"3D",x"87",x"27",x"E1", -- 0x2078
		x"3D",x"87",x"3C",x"87",x"3D",x"87",x"2F",x"0A", -- 0x2080
		x"09",x"02",x"18",x"02",x"15",x"02",x"08",x"02", -- 0x2088
		x"22",x"02",x"23",x"02",x"24",x"02",x"17",x"02", -- 0x2090
		x"18",x"02",x"18",x"02",x"15",x"02",x"2F",x"0A", -- 0x2098
		x"09",x"02",x"18",x"02",x"0B",x"02",x"17",x"02", -- 0x20A0
		x"15",x"02",x"2F",x"0A",x"30",x"0A",x"23",x"02", -- 0x20A8
		x"24",x"02",x"14",x"02",x"2F",x"0A",x"3C",x"02", -- 0x20B0
		x"20",x"E1",x"2E",x"A1",x"31",x"A1",x"22",x"02", -- 0x20B8
		x"11",x"02",x"19",x"02",x"05",x"02",x"0D",x"02", -- 0x20C0
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"02",x"02", -- 0x20C8
		x"22",x"02",x"23",x"02",x"24",x"02",x"22",x"02", -- 0x20D0
		x"23",x"02",x"24",x"02",x"11",x"02",x"10",x"02", -- 0x20D8
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"2F",x"0A", -- 0x20E0
		x"03",x"02",x"19",x"02",x"19",x"02",x"0F",x"02", -- 0x20E8
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"23",x"02", -- 0x20F0
		x"24",x"02",x"0D",x"02",x"32",x"0A",x"24",x"02", -- 0x20F8
		x"25",x"02",x"13",x"02",x"2F",x"0A",x"22",x"02", -- 0x2100
		x"23",x"02",x"24",x"02",x"17",x"02",x"18",x"02", -- 0x2108
		x"15",x"02",x"2F",x"0A",x"30",x"0A",x"23",x"02", -- 0x2110
		x"24",x"02",x"12",x"02",x"31",x"0A",x"25",x"02", -- 0x2118
		x"23",x"02",x"1A",x"02",x"32",x"0A",x"24",x"02", -- 0x2120
		x"22",x"02",x"0C",x"02",x"2F",x"0A",x"22",x"02", -- 0x2128
		x"0E",x"02",x"30",x"0A",x"31",x"0A",x"28",x"42", -- 0x2130
		x"39",x"22",x"39",x"22",x"00",x"00",x"2D",x"42", -- 0x2138
		x"2C",x"22",x"39",x"02",x"00",x"00",x"28",x"42", -- 0x2140
		x"2C",x"42",x"2C",x"22",x"39",x"02",x"2B",x"42", -- 0x2148
		x"2A",x"22",x"2F",x"0A",x"30",x"0A",x"00",x"00", -- 0x2150
		x"00",x"00",x"00",x"00",x"00",x"00",x"2F",x"0A", -- 0x2158
		x"30",x"0A",x"2A",x"42",x"2A",x"22",x"30",x"0A", -- 0x2160
		x"29",x"42",x"2B",x"22",x"31",x"0A",x"32",x"0A", -- 0x2168
		x"2B",x"42",x"2D",x"02",x"2E",x"02",x"2C",x"42", -- 0x2170
		x"2C",x"22",x"39",x"02",x"2C",x"62",x"2A",x"02", -- 0x2178
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"2B",x"62", -- 0x2180
		x"2A",x"02",x"2F",x"0A",x"32",x"0A",x"28",x"62", -- 0x2188
		x"2C",x"62",x"2C",x"02",x"39",x"22",x"2C",x"62", -- 0x2190
		x"2C",x"02",x"2E",x"02",x"00",x"00",x"2F",x"0A", -- 0x2198
		x"2E",x"62",x"39",x"02",x"00",x"00",x"2F",x"0A", -- 0x21A0
		x"09",x"02",x"18",x"02",x"18",x"02",x"22",x"02", -- 0x21A8
		x"24",x"02",x"25",x"02",x"12",x"02",x"23",x"02", -- 0x21B0
		x"22",x"02",x"24",x"02",x"13",x"02",x"24",x"02", -- 0x21B8
		x"25",x"02",x"23",x"02",x"0D",x"02",x"19",x"02", -- 0x21C0
		x"19",x"02",x"0F",x"02",x"2F",x"0A",x"00",x"00", -- 0x21C8
		x"2E",x"62",x"39",x"02",x"39",x"02",x"39",x"62", -- 0x21D0
		x"2C",x"42",x"2A",x"22",x"32",x"0A",x"30",x"0A", -- 0x21D8
		x"31",x"0A",x"09",x"02",x"18",x"02",x"31",x"0A", -- 0x21E0
		x"08",x"02",x"22",x"02",x"23",x"02",x"32",x"0A", -- 0x21E8
		x"09",x"02",x"18",x"02",x"18",x"02",x"0B",x"02", -- 0x21F0
		x"23",x"02",x"24",x"02",x"25",x"02",x"06",x"02", -- 0x21F8
		x"22",x"02",x"23",x"02",x"24",x"02",x"02",x"89", -- 0x2200
		x"09",x"89",x"07",x"89",x"00",x"89",x"3D",x"87", -- 0x2208
		x"3C",x"87",x"3D",x"87",x"19",x"89",x"07",x"89", -- 0x2210
		x"08",x"89",x"05",x"89",x"00",x"00",x"22",x"02", -- 0x2218
		x"11",x"02",x"0F",x"02",x"2F",x"0A",x"2F",x"0A", -- 0x2220
		x"30",x"0A",x"31",x"0A",x"88",x"8C",x"8A",x"8C", -- 0x2228
		x"89",x"8C",x"8B",x"8C",x"8D",x"8C",x"00",x"00", -- 0x2230
		x"88",x"8C",x"89",x"8C",x"5D",x"8C",x"5E",x"8C", -- 0x2238
		x"5F",x"8C",x"85",x"8C",x"8E",x"8C",x"8D",x"8C", -- 0x2240
		x"87",x"8C",x"89",x"8C",x"8B",x"8C",x"40",x"8D", -- 0x2248
		x"6C",x"8C",x"68",x"8C",x"69",x"8C",x"76",x"8C", -- 0x2250
		x"7C",x"8C",x"7D",x"8C",x"89",x"8C",x"8B",x"8C", -- 0x2258
		x"8E",x"8C",x"8F",x"8C",x"8C",x"8C",x"8E",x"8C", -- 0x2260
		x"86",x"8C",x"54",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2268
		x"64",x"8C",x"60",x"8C",x"61",x"8C",x"74",x"8C", -- 0x2270
		x"75",x"8C",x"6D",x"8C",x"78",x"8C",x"79",x"8C", -- 0x2278
		x"89",x"8C",x"8A",x"8C",x"8B",x"8C",x"89",x"8C", -- 0x2280
		x"7A",x"8D",x"7B",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2288
		x"6B",x"8C",x"54",x"8C",x"55",x"8C",x"56",x"8C", -- 0x2290
		x"57",x"8C",x"65",x"8C",x"70",x"8C",x"71",x"8D", -- 0x2298
		x"6F",x"8C",x"5D",x"8C",x"5E",x"8C",x"5F",x"8C", -- 0x22A0
		x"72",x"8C",x"73",x"8C",x"40",x"8D",x"40",x"8D", -- 0x22A8
		x"63",x"8C",x"74",x"8C",x"75",x"8C",x"7C",x"8C", -- 0x22B0
		x"7D",x"8C",x"7A",x"8D",x"7B",x"8C",x"6E",x"8C", -- 0x22B8
		x"67",x"8C",x"74",x"8C",x"75",x"8C",x"50",x"8D", -- 0x22C0
		x"51",x"8D",x"52",x"8D",x"53",x"8D",x"40",x"8D", -- 0x22C8
		x"58",x"8C",x"63",x"8C",x"64",x"8C",x"5B",x"8C", -- 0x22D0
		x"6C",x"8C",x"72",x"8C",x"73",x"8C",x"66",x"8D", -- 0x22D8
		x"50",x"8D",x"53",x"0D",x"52",x"8D",x"53",x"8D", -- 0x22E0
		x"58",x"8C",x"59",x"8C",x"40",x"8D",x"40",x"8D", -- 0x22E8
		x"78",x"8C",x"79",x"8C",x"7E",x"8C",x"7F",x"8C", -- 0x22F0
		x"64",x"8C",x"50",x"8D",x"51",x"8D",x"52",x"8D", -- 0x22F8
		x"53",x"8D",x"76",x"8C",x"6C",x"8C",x"54",x"8C", -- 0x2300
		x"55",x"8C",x"56",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2308
		x"70",x"8C",x"71",x"8D",x"50",x"8D",x"53",x"0D", -- 0x2310
		x"52",x"8D",x"53",x"8D",x"5C",x"8D",x"5D",x"8C", -- 0x2318
		x"5E",x"8C",x"5F",x"8C",x"64",x"8C",x"76",x"8C", -- 0x2320
		x"77",x"8C",x"6D",x"8C",x"40",x"8D",x"67",x"8C", -- 0x2328
		x"72",x"8C",x"7D",x"8C",x"66",x"8D",x"68",x"8C", -- 0x2330
		x"69",x"8C",x"7E",x"8C",x"7F",x"8C",x"7C",x"8C", -- 0x2338
		x"7D",x"8C",x"4C",x"8D",x"4D",x"8D",x"4E",x"8D", -- 0x2340
		x"4F",x"8D",x"65",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2348
		x"55",x"8C",x"56",x"8C",x"57",x"8C",x"60",x"8C", -- 0x2350
		x"61",x"8C",x"6E",x"8C",x"6A",x"8C",x"6B",x"8C", -- 0x2358
		x"77",x"8C",x"44",x"8D",x"45",x"8D",x"46",x"8D", -- 0x2360
		x"47",x"8D",x"74",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2368
		x"6B",x"8C",x"58",x"8C",x"59",x"8C",x"5A",x"8C", -- 0x2370
		x"5B",x"8C",x"66",x"8D",x"62",x"8C",x"63",x"8C", -- 0x2378
		x"6A",x"8C",x"6B",x"8C",x"5C",x"8D",x"5D",x"8C", -- 0x2380
		x"5E",x"8C",x"5F",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2388
		x"63",x"8C",x"74",x"8C",x"75",x"8C",x"78",x"8C", -- 0x2390
		x"79",x"8C",x"7E",x"8C",x"7F",x"8C",x"6F",x"8C", -- 0x2398
		x"62",x"8C",x"63",x"8C",x"7C",x"8C",x"7D",x"8C", -- 0x23A0
		x"77",x"8C",x"69",x"8C",x"40",x"8D",x"40",x"8D", -- 0x23A8
		x"49",x"8D",x"4A",x"8D",x"4B",x"8D",x"78",x"8C", -- 0x23B0
		x"79",x"8C",x"7E",x"8C",x"7F",x"8C",x"67",x"8C", -- 0x23B8
		x"76",x"8C",x"54",x"8C",x"55",x"8C",x"56",x"8C", -- 0x23C0
		x"57",x"8C",x"61",x"8C",x"40",x"8D",x"40",x"8D", -- 0x23C8
		x"41",x"8D",x"42",x"8D",x"43",x"8D",x"70",x"8C", -- 0x23D0
		x"71",x"8D",x"77",x"8C",x"54",x"8C",x"55",x"8C", -- 0x23D8
		x"56",x"8C",x"57",x"8C",x"6C",x"8C",x"77",x"8C", -- 0x23E0
		x"6A",x"8C",x"6B",x"8C",x"40",x"8D",x"76",x"8C", -- 0x23E8
		x"7A",x"8D",x"7B",x"8C",x"7C",x"8C",x"7D",x"8C", -- 0x23F0
		x"58",x"8C",x"59",x"8C",x"5A",x"8C",x"5B",x"8C", -- 0x23F8
		x"7E",x"8C",x"7F",x"8C",x"64",x"8C",x"6F",x"8C", -- 0x2400
		x"62",x"8C",x"63",x"8C",x"40",x"8D",x"5F",x"8C", -- 0x2408
		x"72",x"8C",x"73",x"8C",x"54",x"8C",x"55",x"8C", -- 0x2410
		x"56",x"8C",x"57",x"8C",x"6D",x"8C",x"9C",x"86", -- 0x2418
		x"9D",x"86",x"9E",x"86",x"9F",x"86",x"67",x"8C", -- 0x2420
		x"58",x"8C",x"59",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2428
		x"5F",x"8C",x"68",x"8C",x"69",x"8C",x"74",x"8C", -- 0x2430
		x"75",x"8C",x"6C",x"8C",x"65",x"8C",x"94",x"86", -- 0x2438
		x"95",x"86",x"96",x"86",x"97",x"86",x"7A",x"8D", -- 0x2440
		x"7B",x"8C",x"77",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2448
		x"57",x"8C",x"60",x"8C",x"61",x"8C",x"6F",x"8C", -- 0x2450
		x"76",x"8C",x"64",x"8C",x"6E",x"8C",x"98",x"86", -- 0x2458
		x"99",x"86",x"9A",x"86",x"9B",x"86",x"72",x"8C", -- 0x2460
		x"73",x"8C",x"78",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2468
		x"5E",x"8C",x"5F",x"8C",x"6D",x"8C",x"90",x"86", -- 0x2470
		x"91",x"86",x"92",x"86",x"93",x"86",x"6C",x"8C", -- 0x2478
		x"6D",x"8C",x"70",x"8C",x"40",x"8D",x"40",x"8D", -- 0x2480
		x"7E",x"8C",x"7F",x"8C",x"65",x"8C",x"74",x"8C", -- 0x2488
		x"75",x"8C",x"82",x"8C",x"83",x"8C",x"7E",x"8C", -- 0x2490
		x"7F",x"8C",x"6A",x"8C",x"6B",x"8C",x"64",x"8C", -- 0x2498
		x"65",x"8C",x"6E",x"8C",x"40",x"8D",x"40",x"8D", -- 0x24A0
		x"55",x"8C",x"56",x"8C",x"57",x"8C",x"82",x"8C", -- 0x24A8
		x"85",x"8C",x"8E",x"8C",x"8C",x"8C",x"86",x"8C", -- 0x24B0
		x"76",x"8C",x"62",x"8C",x"63",x"8C",x"68",x"8C", -- 0x24B8
		x"69",x"8C",x"66",x"8D",x"40",x"8D",x"40",x"8D", -- 0x24C0
		x"82",x"8C",x"83",x"8C",x"81",x"8C",x"87",x"8C", -- 0x24C8
		x"83",x"8C",x"7C",x"8C",x"7D",x"8C",x"60",x"8C", -- 0x24D0
		x"61",x"8C",x"74",x"8C",x"40",x"8D",x"8C",x"8C", -- 0x24D8
		x"8E",x"8C",x"80",x"8C",x"81",x"8C",x"82",x"8C", -- 0x24E0
		x"83",x"8C",x"81",x"8C",x"40",x"8D",x"8E",x"8C", -- 0x24E8
		x"8F",x"8C",x"8D",x"8C",x"8C",x"8C",x"40",x"8D", -- 0x24F0
		x"8E",x"8C",x"8F",x"8C",x"8D",x"8C",x"2F",x"0A", -- 0x24F8
		x"8D",x"8C",x"30",x"0A",x"8D",x"8C",x"31",x"0A", -- 0x2500
		x"8C",x"8C",x"8F",x"8C",x"8E",x"8C",x"8C",x"8C", -- 0x2508
		x"8F",x"8C",x"8E",x"8C",x"31",x"0A",x"30",x"0A", -- 0x2510
		x"31",x"0A",x"32",x"0A",x"8D",x"8C",x"8F",x"8C", -- 0x2518
		x"8D",x"8C",x"2F",x"03",x"8C",x"8C",x"89",x"8C", -- 0x2520
		x"5D",x"8C",x"5E",x"8C",x"5F",x"8C",x"5E",x"8C", -- 0x2528
		x"5F",x"8C",x"76",x"8C",x"5D",x"8C",x"85",x"8C", -- 0x2530
		x"8C",x"8C",x"8F",x"8C",x"8D",x"8C",x"66",x"8D", -- 0x2538
		x"5D",x"8C",x"5E",x"8C",x"5F",x"8C",x"56",x"07", -- 0x2540
		x"5E",x"07",x"57",x"07",x"5E",x"07",x"5E",x"07", -- 0x2548
		x"3C",x"87",x"3D",x"87",x"3C",x"87",x"5A",x"07", -- 0x2550
		x"59",x"07",x"5A",x"07",x"5B",x"07",x"5A",x"07", -- 0x2558
		x"5F",x"07",x"5E",x"07",x"58",x"07",x"56",x"07", -- 0x2560
		x"5E",x"07",x"58",x"07",x"40",x"07",x"59",x"07", -- 0x2568
		x"5B",x"07",x"59",x"07",x"5A",x"07",x"59",x"07", -- 0x2570
		x"5A",x"07",x"5C",x"07",x"5B",x"07",x"5D",x"07", -- 0x2578
		x"3C",x"87",x"3D",x"87",x"3C",x"87",x"40",x"07", -- 0x2580
		x"55",x"07",x"5E",x"07",x"5B",x"07",x"5C",x"07", -- 0x2588
		x"5B",x"07",x"59",x"07",x"5A",x"07",x"5F",x"07", -- 0x2590
		x"54",x"07",x"5E",x"07",x"5E",x"07",x"5B",x"07", -- 0x2598
		x"5A",x"07",x"5B",x"07",x"59",x"07",x"88",x"8C", -- 0x25A0
		x"8B",x"8C",x"59",x"07",x"5A",x"07",x"66",x"8D", -- 0x25A8
		x"5D",x"8C",x"5E",x"8C",x"55",x"8C",x"40",x"07", -- 0x25B0
		x"80",x"8C",x"82",x"8C",x"76",x"8C",x"40",x"07", -- 0x25B8
		x"8C",x"8C",x"8E",x"8C",x"86",x"8C",x"40",x"07", -- 0x25C0
		x"31",x"0A",x"8F",x"8C",x"80",x"8C",x"83",x"8C", -- 0x25C8
		x"76",x"8C",x"64",x"8C",x"77",x"8C",x"40",x"07", -- 0x25D0
		x"32",x"0A",x"8D",x"8C",x"8C",x"8C",x"8E",x"8C", -- 0x25D8
		x"86",x"8C",x"74",x"8C",x"75",x"8C",x"81",x"8C", -- 0x25E0
		x"8D",x"8C",x"8C",x"8C",x"80",x"8C",x"8F",x"8C", -- 0x25E8
		x"80",x"8C",x"83",x"8C",x"82",x"8C",x"8D",x"8C", -- 0x25F0
		x"8C",x"8C",x"2F",x"0A",x"8F",x"8C",x"33",x"02", -- 0x25F8
		x"2F",x"0A",x"34",x"02",x"30",x"0A",x"31",x"0A", -- 0x2600
		x"33",x"02",x"32",x"0A",x"33",x"02",x"33",x"02", -- 0x2608
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"2F",x"0A", -- 0x2610
		x"34",x"02",x"32",x"0A",x"30",x"0A",x"31",x"0A", -- 0x2618
		x"33",x"02",x"34",x"02",x"32",x"0A",x"2F",x"0A", -- 0x2620
		x"30",x"0A",x"33",x"02",x"34",x"02",x"35",x"02", -- 0x2628
		x"3C",x"02",x"3D",x"02",x"3B",x"02",x"3B",x"02", -- 0x2630
		x"3D",x"02",x"35",x"02",x"3C",x"02",x"3C",x"02", -- 0x2638
		x"3B",x"02",x"35",x"02",x"3D",x"02",x"36",x"02", -- 0x2640
		x"3C",x"02",x"35",x"02",x"3B",x"02",x"3C",x"02", -- 0x2648
		x"36",x"02",x"3B",x"02",x"3D",x"02",x"36",x"02", -- 0x2650
		x"35",x"02",x"35",x"02",x"36",x"02",x"3B",x"02", -- 0x2658
		x"3C",x"02",x"3D",x"02",x"35",x"02",x"31",x"E1", -- 0x2660
		x"27",x"C1",x"3C",x"87",x"3D",x"87",x"38",x"81", -- 0x2668
		x"20",x"A1",x"3B",x"02",x"3C",x"02",x"3C",x"87", -- 0x2670
		x"25",x"81",x"3C",x"02",x"3D",x"02",x"3D",x"87", -- 0x2678
		x"3C",x"87",x"21",x"A1",x"3C",x"02",x"3C",x"87", -- 0x2680
		x"3D",x"87",x"27",x"81",x"31",x"A1",x"2F",x"0A", -- 0x2688
		x"30",x"0A",x"2B",x"62",x"3B",x"02",x"30",x"0A", -- 0x2690
		x"31",x"0A",x"29",x"62",x"3C",x"02",x"2D",x"62", -- 0x2698
		x"3B",x"02",x"3C",x"02",x"3D",x"02",x"38",x"42", -- 0x26A0
		x"3D",x"02",x"3B",x"02",x"3C",x"02",x"29",x"62", -- 0x26A8
		x"3C",x"02",x"3D",x"02",x"3B",x"02",x"2F",x"0A", -- 0x26B0
		x"2E",x"62",x"39",x"02",x"00",x"02",x"15",x"02", -- 0x26B8
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"23",x"02", -- 0x26C0
		x"14",x"02",x"2F",x"0A",x"32",x"0A",x"22",x"02", -- 0x26C8
		x"23",x"02",x"24",x"02",x"1A",x"02",x"14",x"02", -- 0x26D0
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"24",x"02", -- 0x26D8
		x"17",x"02",x"15",x"02",x"2F",x"0A",x"25",x"02", -- 0x26E0
		x"24",x"02",x"23",x"02",x"1A",x"02",x"23",x"02", -- 0x26E8
		x"11",x"02",x"0F",x"02",x"30",x"0A",x"0E",x"02", -- 0x26F0
		x"30",x"0A",x"31",x"0A",x"32",x"0A",x"24",x"02", -- 0x26F8
		x"25",x"02",x"23",x"02",x"1A",x"02",x"22",x"02", -- 0x2700
		x"23",x"02",x"0E",x"02",x"2F",x"0A",x"19",x"02", -- 0x2708
		x"0F",x"02",x"2F",x"0A",x"30",x"0A",x"44",x"23", -- 0x2710
		x"4E",x"23",x"4E",x"63",x"41",x"63",x"40",x"63", -- 0x2718
		x"42",x"63",x"44",x"63",x"40",x"03",x"4A",x"03", -- 0x2720
		x"49",x"43",x"43",x"43",x"2F",x"0A",x"2F",x"0A", -- 0x2728
		x"41",x"03",x"4E",x"03",x"51",x"03",x"4E",x"43", -- 0x2730
		x"41",x"43",x"41",x"23",x"40",x"03",x"30",x"0A", -- 0x2738
		x"44",x"23",x"4E",x"23",x"51",x"23",x"51",x"23", -- 0x2740
		x"4E",x"63",x"41",x"63",x"30",x"0A",x"2F",x"0A", -- 0x2748
		x"45",x"03",x"4A",x"03",x"4B",x"03",x"44",x"63", -- 0x2750
		x"45",x"03",x"4B",x"03",x"40",x"03",x"31",x"0A", -- 0x2758
		x"44",x"03",x"42",x"03",x"47",x"03",x"45",x"43", -- 0x2760
		x"44",x"03",x"40",x"03",x"40",x"03",x"48",x"03", -- 0x2768
		x"49",x"03",x"4A",x"03",x"4B",x"03",x"44",x"63", -- 0x2770
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"1B",x"02", -- 0x2778
		x"22",x"02",x"23",x"02",x"24",x"02",x"04",x"02", -- 0x2780
		x"05",x"02",x"25",x"02",x"22",x"02",x"2F",x"0A", -- 0x2788
		x"30",x"0A",x"01",x"02",x"23",x"02",x"30",x"0A", -- 0x2790
		x"31",x"0A",x"1B",x"02",x"25",x"02",x"31",x"0A", -- 0x2798
		x"32",x"0A",x"00",x"02",x"24",x"02",x"32",x"0A", -- 0x27A0
		x"2F",x"0A",x"30",x"0A",x"01",x"02",x"2F",x"0A", -- 0x27A8
		x"30",x"0A",x"31",x"0A",x"04",x"02",x"05",x"02", -- 0x27B0
		x"23",x"02",x"24",x"02",x"25",x"02",x"09",x"02", -- 0x27B8
		x"18",x"02",x"18",x"02",x"16",x"02",x"22",x"02", -- 0x27C0
		x"24",x"02",x"25",x"02",x"13",x"02",x"2F",x"0A", -- 0x27C8
		x"02",x"02",x"23",x"02",x"24",x"02",x"30",x"0A", -- 0x27D0
		x"31",x"0A",x"32",x"0A",x"03",x"02",x"40",x"03", -- 0x27D8
		x"42",x"03",x"42",x"03",x"40",x"03",x"4F",x"63", -- 0x27E0
		x"4E",x"63",x"42",x"23",x"44",x"63",x"41",x"03", -- 0x27E8
		x"4E",x"03",x"4F",x"03",x"46",x"63",x"2F",x"0A", -- 0x27F0
		x"30",x"0A",x"31",x"0A",x"46",x"03",x"48",x"63", -- 0x27F8
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"31",x"0A", -- 0x2800
		x"32",x"0A",x"2F",x"0A",x"44",x"03",x"47",x"03", -- 0x2808
		x"43",x"63",x"2F",x"0A",x"32",x"0A",x"45",x"03", -- 0x2810
		x"45",x"43",x"31",x"0A",x"30",x"0A",x"46",x"23", -- 0x2818
		x"45",x"43",x"2F",x"0A",x"32",x"0A",x"2F",x"0A", -- 0x2820
		x"30",x"0A",x"31",x"0A",x"48",x"23",x"49",x"43", -- 0x2828
		x"43",x"43",x"32",x"0A",x"2F",x"0A",x"31",x"0A", -- 0x2830
		x"32",x"0A",x"43",x"23",x"49",x"43",x"2F",x"0A", -- 0x2838
		x"30",x"0A",x"46",x"23",x"45",x"43",x"32",x"0A", -- 0x2840
		x"43",x"23",x"49",x"43",x"43",x"43",x"30",x"0A", -- 0x2848
		x"45",x"03",x"46",x"43",x"32",x"0A",x"31",x"0A", -- 0x2850
		x"2F",x"0A",x"48",x"03",x"46",x"63",x"43",x"63", -- 0x2858
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"2F",x"0A", -- 0x2860
		x"30",x"0A",x"31",x"0A",x"43",x"03",x"46",x"63", -- 0x2868
		x"31",x"0A",x"32",x"0A",x"2F",x"0A",x"46",x"03", -- 0x2870
		x"43",x"63",x"2F",x"0A",x"30",x"0A",x"43",x"23", -- 0x2878
		x"4A",x"03",x"45",x"43",x"2F",x"0A",x"45",x"03", -- 0x2880
		x"49",x"03",x"43",x"43",x"32",x"0A",x"46",x"23", -- 0x2888
		x"48",x"43",x"30",x"0A",x"9C",x"02",x"46",x"43", -- 0x2890
		x"96",x"02",x"97",x"02",x"98",x"02",x"43",x"43", -- 0x2898
		x"90",x"02",x"91",x"02",x"92",x"02",x"2F",x"0A", -- 0x28A0
		x"30",x"0A",x"45",x"03",x"45",x"43",x"30",x"0A", -- 0x28A8
		x"31",x"0A",x"43",x"03",x"47",x"63",x"BC",x"02", -- 0x28B0
		x"2F",x"0A",x"30",x"0A",x"48",x"03",x"47",x"63", -- 0x28B8
		x"41",x"63",x"2F",x"0A",x"30",x"0A",x"41",x"03", -- 0x28C0
		x"47",x"03",x"40",x"63",x"42",x"23",x"42",x"23", -- 0x28C8
		x"40",x"23",x"40",x"43",x"40",x"03",x"2F",x"0A", -- 0x28D0
		x"45",x"03",x"47",x"43",x"42",x"03",x"30",x"0A", -- 0x28D8
		x"45",x"03",x"45",x"43",x"31",x"0A",x"31",x"0A", -- 0x28E0
		x"43",x"03",x"46",x"63",x"32",x"0A",x"2F",x"0A", -- 0x28E8
		x"30",x"0A",x"46",x"03",x"43",x"63",x"31",x"0A", -- 0x28F0
		x"32",x"0A",x"43",x"03",x"47",x"63",x"30",x"0A", -- 0x28F8
		x"31",x"0A",x"32",x"0A",x"48",x"03",x"43",x"03", -- 0x2900
		x"47",x"63",x"42",x"23",x"40",x"03",x"32",x"0A", -- 0x2908
		x"41",x"03",x"42",x"03",x"40",x"03",x"22",x"02", -- 0x2910
		x"23",x"02",x"17",x"02",x"15",x"02",x"80",x"02", -- 0x2918
		x"BA",x"02",x"BB",x"02",x"BC",x"02",x"80",x"02", -- 0x2920
		x"B3",x"02",x"B4",x"02",x"B5",x"02",x"B6",x"02", -- 0x2928
		x"2F",x"0A",x"30",x"0A",x"31",x"0A",x"00",x"00", -- 0x2930
		x"AC",x"02",x"AD",x"02",x"AE",x"02",x"AF",x"02", -- 0x2938
		x"30",x"0A",x"31",x"0A",x"32",x"0A",x"00",x"00", -- 0x2940
		x"A6",x"02",x"A7",x"02",x"A8",x"02",x"2F",x"0A", -- 0x2948
		x"30",x"0A",x"31",x"0A",x"9C",x"02",x"00",x"00", -- 0x2950
		x"00",x"00",x"00",x"00",x"00",x"00",x"9D",x"02", -- 0x2958
		x"9E",x"02",x"9F",x"02",x"80",x"02",x"2F",x"0A", -- 0x2960
		x"96",x"02",x"97",x"02",x"98",x"02",x"99",x"02", -- 0x2968
		x"9A",x"02",x"9B",x"02",x"80",x"02",x"30",x"0A", -- 0x2970
		x"90",x"02",x"91",x"02",x"92",x"02",x"93",x"02", -- 0x2978
		x"94",x"02",x"95",x"02",x"80",x"02",x"89",x"02", -- 0x2980
		x"8A",x"02",x"8B",x"02",x"8C",x"02",x"8D",x"02", -- 0x2988
		x"8E",x"02",x"8F",x"02",x"90",x"02",x"2F",x"0A", -- 0x2990
		x"83",x"02",x"84",x"02",x"85",x"02",x"86",x"02", -- 0x2998
		x"87",x"02",x"88",x"02",x"80",x"02",x"80",x"02", -- 0x29A0
		x"81",x"02",x"82",x"02",x"80",x"02",x"9F",x"02", -- 0x29A8
		x"BD",x"02",x"BE",x"02",x"BF",x"02",x"9B",x"02", -- 0x29B0
		x"B7",x"02",x"B8",x"02",x"B9",x"02",x"BA",x"02", -- 0x29B8
		x"BB",x"02",x"BC",x"02",x"2F",x"0A",x"95",x"02", -- 0x29C0
		x"B0",x"02",x"B1",x"02",x"B2",x"02",x"B3",x"02", -- 0x29C8
		x"B4",x"02",x"B5",x"02",x"B6",x"02",x"8F",x"02", -- 0x29D0
		x"A9",x"02",x"AA",x"02",x"AB",x"02",x"AC",x"02", -- 0x29D8
		x"AD",x"02",x"AE",x"02",x"AF",x"02",x"88",x"02", -- 0x29E0
		x"A3",x"02",x"A4",x"02",x"A5",x"02",x"A6",x"02", -- 0x29E8
		x"A7",x"02",x"A8",x"02",x"30",x"0A",x"82",x"02", -- 0x29F0
		x"A0",x"02",x"A1",x"02",x"A2",x"02",x"80",x"02", -- 0x29F8
		x"BF",x"02",x"2F",x"0A",x"30",x"0A",x"80",x"02", -- 0x2A00
		x"B9",x"02",x"BA",x"02",x"BB",x"02",x"80",x"02", -- 0x2A08
		x"B2",x"02",x"B3",x"02",x"B4",x"02",x"B5",x"02", -- 0x2A10
		x"B6",x"02",x"31",x"0A",x"32",x"0A",x"80",x"02", -- 0x2A18
		x"AB",x"02",x"AC",x"02",x"AD",x"02",x"AE",x"02", -- 0x2A20
		x"AF",x"02",x"30",x"0A",x"31",x"0A",x"80",x"02", -- 0x2A28
		x"A5",x"02",x"A6",x"02",x"A7",x"02",x"A8",x"02", -- 0x2A30
		x"30",x"0A",x"31",x"0A",x"32",x"0A",x"80",x"02", -- 0x2A38
		x"A2",x"02",x"30",x"0A",x"2F",x"0A",x"2F",x"0A", -- 0x2A40
		x"9C",x"02",x"9D",x"02",x"9E",x"02",x"97",x"02", -- 0x2A48
		x"98",x"02",x"99",x"02",x"9A",x"02",x"91",x"02", -- 0x2A50
		x"92",x"02",x"93",x"02",x"94",x"02",x"8B",x"02", -- 0x2A58
		x"8C",x"02",x"8D",x"02",x"8E",x"02",x"84",x"02", -- 0x2A60
		x"85",x"02",x"86",x"02",x"87",x"02",x"2F",x"0A", -- 0x2A68
		x"30",x"0A",x"80",x"02",x"81",x"02",x"2F",x"0A", -- 0x2A70
		x"30",x"0A",x"31",x"0A",x"96",x"02",x"32",x"0A", -- 0x2A78
		x"2F",x"0A",x"30",x"0A",x"90",x"02",x"31",x"0A", -- 0x2A80
		x"32",x"0A",x"89",x"02",x"8A",x"02",x"2F",x"0A", -- 0x2A88
		x"30",x"0A",x"32",x"0A",x"83",x"02",x"22",x"02", -- 0x2A90
		x"23",x"02",x"17",x"02",x"00",x"02",x"01",x"02", -- 0x2A98
		x"22",x"02",x"23",x"02",x"24",x"02",x"00",x"02", -- 0x2AA0
		x"23",x"02",x"24",x"02",x"25",x"02",x"02",x"02", -- 0x2AA8
		x"19",x"02",x"19",x"02",x"10",x"02",x"05",x"02", -- 0x2AB0
		x"22",x"02",x"23",x"02",x"00",x"02",x"1B",x"02", -- 0x2AB8
		x"23",x"02",x"24",x"02",x"25",x"02",x"FD",x"03", -- 0x2AC0
		x"FD",x"03",x"FD",x"03",x"FD",x"03",x"4A",x"03", -- 0x2AC8
		x"4B",x"03",x"4A",x"03",x"4B",x"03",x"4B",x"03", -- 0x2AD0
		x"4A",x"03",x"4B",x"03",x"4A",x"03",x"39",x"22", -- 0x2AD8
		x"2C",x"42",x"2C",x"22",x"39",x"02",x"1B",x"02", -- 0x2AE0
		x"22",x"02",x"23",x"02",x"24",x"02",x"1C",x"89", -- 0x2AE8
		x"11",x"C9",x"3C",x"87",x"3D",x"87",x"3C",x"02", -- 0x2AF0
		x"3D",x"02",x"20",x"C1",x"31",x"81",x"2F",x"0A", -- 0x2AF8
		x"30",x"0A",x"2E",x"62",x"00",x"00",x"22",x"02", -- 0x2B00
		x"23",x"02",x"24",x"02",x"0C",x"02",x"09",x"02", -- 0x2B08
		x"18",x"02",x"18",x"02",x"00",x"00",x"2F",x"0A", -- 0x2B10
		x"30",x"0A",x"02",x"02",x"23",x"02",x"3C",x"02", -- 0x2B18
		x"3D",x"02",x"20",x"E1",x"38",x"C1",x"3C",x"87", -- 0x2B20
		x"BE",x"8E",x"B7",x"8E",x"B7",x"8E",x"B7",x"8E", -- 0x2B28
		x"B7",x"8E",x"BF",x"8E",x"79",x"0E",x"3D",x"87", -- 0x2B30
		x"BD",x"8E",x"EC",x"00",x"BC",x"8E",x"BC",x"CE", -- 0x2B38
		x"74",x"00",x"C1",x"8E",x"7A",x"0E",x"3C",x"87", -- 0x2B40
		x"B5",x"8E",x"E4",x"00",x"BC",x"8E",x"BC",x"CE", -- 0x2B48
		x"73",x"00",x"C0",x"8E",x"AF",x"8E",x"AC",x"8F", -- 0x2B50
		x"AD",x"8E",x"FF",x"00",x"AE",x"8E",x"AE",x"CE", -- 0x2B58
		x"DE",x"00",x"AD",x"CE",x"CF",x"8B",x"A4",x"8F", -- 0x2B60
		x"A5",x"8E",x"D7",x"80",x"BC",x"8E",x"BC",x"CE", -- 0x2B68
		x"74",x"00",x"A5",x"CE",x"C7",x"8B",x"B8",x"8E", -- 0x2B70
		x"BB",x"8E",x"EC",x"00",x"BC",x"8E",x"BC",x"CE", -- 0x2B78
		x"73",x"00",x"DF",x"00",x"C3",x"8E",x"B0",x"8E", -- 0x2B80
		x"A3",x"80",x"E4",x"00",x"BC",x"8E",x"BC",x"CE", -- 0x2B88
		x"ED",x"00",x"EE",x"00",x"EF",x"00",x"A8",x"8E", -- 0x2B90
		x"BB",x"8E",x"EC",x"00",x"BC",x"8E",x"E0",x"0E", -- 0x2B98
		x"E5",x"00",x"E6",x"00",x"E7",x"00",x"A0",x"8E", -- 0x2BA0
		x"A3",x"80",x"E4",x"00",x"BC",x"8E",x"F0",x"0E", -- 0x2BA8
		x"F1",x"00",x"F2",x"00",x"FE",x"00",x"7A",x"0E", -- 0x2BB0
		x"75",x"2E",x"3C",x"87",x"3D",x"87",x"B9",x"8E", -- 0x2BB8
		x"AA",x"8E",x"FF",x"00",x"AE",x"8E",x"E8",x"0E", -- 0x2BC0
		x"E9",x"00",x"EA",x"00",x"EB",x"00",x"7A",x"0E", -- 0x2BC8
		x"76",x"2E",x"3D",x"87",x"3D",x"87",x"B1",x"8E", -- 0x2BD0
		x"BB",x"8E",x"EC",x"00",x"A2",x"8E",x"BC",x"CE", -- 0x2BD8
		x"E1",x"00",x"E2",x"00",x"E3",x"00",x"7A",x"0E", -- 0x2BE0
		x"77",x"2E",x"3D",x"87",x"3C",x"87",x"A9",x"8E", -- 0x2BE8
		x"A3",x"80",x"E4",x"00",x"A2",x"8E",x"BC",x"CE", -- 0x2BF0
		x"DC",x"80",x"DD",x"80",x"DE",x"8B",x"79",x"2E", -- 0x2BF8
		x"78",x"0E",x"3D",x"87",x"3C",x"87",x"A1",x"8E", -- 0x2C00
		x"BB",x"8E",x"EC",x"00",x"A2",x"8E",x"BC",x"CE", -- 0x2C08
		x"D4",x"80",x"D5",x"80",x"D6",x"8B",x"BA",x"8E", -- 0x2C10
		x"A3",x"80",x"E4",x"00",x"A2",x"8E",x"BC",x"CE", -- 0x2C18
		x"CC",x"80",x"CD",x"80",x"CE",x"8B",x"3C",x"87", -- 0x2C20
		x"B3",x"8E",x"FF",x"00",x"AE",x"8E",x"AE",x"CE", -- 0x2C28
		x"C4",x"8E",x"C5",x"80",x"7A",x"0E",x"3D",x"87", -- 0x2C30
		x"AB",x"8E",x"D7",x"80",x"BC",x"8E",x"BC",x"CE", -- 0x2C38
		x"DF",x"00",x"C2",x"8E",x"79",x"2E",x"3C",x"87", -- 0x2C40
		x"D8",x"8E",x"D9",x"8E",x"DA",x"8E",x"DA",x"CE", -- 0x2C48
		x"D9",x"CE",x"DB",x"8E",x"7B",x"0E",x"3D",x"87", -- 0x2C50
		x"D0",x"8E",x"D1",x"8E",x"D2",x"8E",x"D2",x"CE", -- 0x2C58
		x"D1",x"CE",x"D3",x"8E",x"7E",x"2E",x"3C",x"87", -- 0x2C60
		x"C8",x"8E",x"C9",x"8E",x"CA",x"8E",x"CA",x"CE", -- 0x2C68
		x"C9",x"CE",x"CB",x"8E",x"3D",x"87",x"3D",x"87", -- 0x2C70
		x"3C",x"87",x"A6",x"8B",x"A7",x"8B",x"A7",x"CB", -- 0x2C78
		x"A6",x"CB",x"3D",x"87",x"3C",x"87",x"3C",x"87", -- 0x2C80
		x"7E",x"4E",x"7C",x"0E",x"7C",x"0E",x"7C",x"0E", -- 0x2C88
		x"7C",x"0E",x"7C",x"0E",x"7F",x"0E",x"77",x"0E", -- 0x2C90
		x"3C",x"87",x"3D",x"87",x"3C",x"8E",x"76",x"0E", -- 0x2C98
		x"3C",x"87",x"3D",x"C7",x"3C",x"87",x"75",x"0E", -- 0x2CA0
		x"3C",x"87",x"3D",x"87",x"3C",x"8E",x"79",x"0E", -- 0x2CA8
		x"78",x"0E",x"3C",x"87",x"3D",x"87",x"7A",x"0E", -- 0x2CB0
		x"77",x"0E",x"3D",x"87",x"3C",x"87",x"7A",x"0E", -- 0x2CB8
		x"76",x"0E",x"3C",x"87",x"3D",x"87",x"7A",x"0E", -- 0x2CC0
		x"75",x"0E",x"3D",x"87",x"3C",x"87",x"77",x"2E", -- 0x2CC8
		x"3C",x"87",x"3D",x"87",x"3C",x"87",x"7D",x"2E", -- 0x2CD0
		x"3C",x"87",x"3D",x"87",x"3C",x"87",x"75",x"2E", -- 0x2CD8
		x"3D",x"87",x"3C",x"87",x"3D",x"87",x"78",x"2E", -- 0x2CE0
		x"3D",x"87",x"3C",x"87",x"3D",x"87",x"00",x"89", -- 0x2CE8
		x"22",x"02",x"23",x"02",x"17",x"02",x"22",x"02", -- 0x2CF0
		x"11",x"02",x"19",x"02",x"19",x"02",x"31",x"00", -- 0x2CF8
		x"F0",x"21",x"00",x"D0",x"CD",x"82",x"AD",x"21", -- 0x2D00
		x"00",x"D8",x"11",x"00",x"04",x"CD",x"85",x"AD", -- 0x2D08
		x"21",x"00",x"E0",x"CD",x"82",x"AD",x"31",x"00", -- 0x2D10
		x"E8",x"21",x"00",x"E8",x"CD",x"82",x"AD",x"CD", -- 0x2D18
		x"03",x"AF",x"16",x"3C",x"01",x"08",x"10",x"21", -- 0x2D20
		x"AD",x"D5",x"CD",x"53",x"02",x"16",x"3D",x"01", -- 0x2D28
		x"02",x"10",x"21",x"AD",x"D5",x"CD",x"53",x"02", -- 0x2D30
		x"21",x"50",x"B8",x"CD",x"22",x"02",x"21",x"34", -- 0x2D38
		x"D3",x"11",x"40",x"B8",x"CD",x"26",x"AE",x"DD", -- 0x2D40
		x"21",x"00",x"E0",x"FD",x"21",x"B4",x"D1",x"CD", -- 0x2D48
		x"C6",x"AD",x"DD",x"21",x"00",x"E8",x"CD",x"C6", -- 0x2D50
		x"AD",x"DD",x"21",x"00",x"D0",x"CD",x"C6",x"AD", -- 0x2D58
		x"DD",x"21",x"00",x"D8",x"CD",x"C6",x"AD",x"CD", -- 0x2D60
		x"E0",x"11",x"21",x"00",x"E0",x"11",x"01",x"E0", -- 0x2D68
		x"01",x"FF",x"0F",x"36",x"00",x"ED",x"B0",x"CD", -- 0x2D70
		x"16",x"04",x"01",x"3B",x"AE",x"AF",x"FF",x"C3", -- 0x2D78
		x"84",x"00",x"11",x"00",x"08",x"06",x"01",x"D5", -- 0x2D80
		x"E5",x"48",x"71",x"CB",x"01",x"23",x"1B",x"7A", -- 0x2D88
		x"B3",x"20",x"F7",x"E1",x"D1",x"48",x"D5",x"E5", -- 0x2D90
		x"79",x"BE",x"20",x"1A",x"CB",x"01",x"23",x"1B", -- 0x2D98
		x"7A",x"B3",x"20",x"F4",x"E1",x"D1",x"CB",x"00", -- 0x2DA0
		x"30",x"DD",x"06",x"04",x"36",x"00",x"23",x"10", -- 0x2DA8
		x"FB",x"C9",x"06",x"07",x"18",x"F6",x"DD",x"E1", -- 0x2DB0
		x"D1",x"DD",x"75",x"00",x"DD",x"74",x"01",x"DD", -- 0x2DB8
		x"71",x"02",x"DD",x"77",x"03",x"C9",x"FD",x"E5", -- 0x2DC0
		x"E1",x"DD",x"7E",x"01",x"DD",x"BE",x"00",x"28", -- 0x2DC8
		x"28",x"CD",x"06",x"AE",x"DD",x"7E",x"00",x"CD", -- 0x2DD0
		x"06",x"AE",x"09",x"DD",x"7E",x"02",x"CD",x"06", -- 0x2DD8
		x"AE",x"09",x"DD",x"7E",x"03",x"CD",x"06",x"AE", -- 0x2DE0
		x"FD",x"E5",x"E1",x"01",x"00",x"04",x"09",x"16", -- 0x2DE8
		x"16",x"01",x"01",x"11",x"CD",x"53",x"02",x"18", -- 0x2DF0
		x"08",x"11",x"28",x"B8",x"06",x"0A",x"CD",x"EE", -- 0x2DF8
		x"01",x"FD",x"2B",x"FD",x"2B",x"C9",x"F5",x"0F", -- 0x2E00
		x"0F",x"0F",x"0F",x"CD",x"0F",x"AE",x"F1",x"E6", -- 0x2E08
		x"0F",x"77",x"01",x"20",x"00",x"09",x"C9",x"C5", -- 0x2E10
		x"D5",x"E5",x"CD",x"EE",x"01",x"E1",x"2B",x"2B", -- 0x2E18
		x"D1",x"C1",x"0D",x"20",x"F2",x"C9",x"1A",x"B7", -- 0x2E20
		x"C8",x"13",x"E5",x"47",x"CD",x"EE",x"01",x"E1", -- 0x2E28
		x"2B",x"2B",x"18",x"F2",x"71",x"0C",x"2B",x"2B", -- 0x2E30
		x"10",x"FA",x"C9",x"CD",x"85",x"02",x"3E",x"02", -- 0x2E38
		x"32",x"3A",x"EC",x"CD",x"A7",x"02",x"CD",x"24", -- 0x2E40
		x"B7",x"CD",x"75",x"B7",x"06",x"02",x"DF",x"3A", -- 0x2E48
		x"01",x"C0",x"2F",x"E6",x"0F",x"28",x"F5",x"06", -- 0x2E50
		x"02",x"DF",x"3A",x"01",x"C0",x"2F",x"E6",x"0F", -- 0x2E58
		x"20",x"F5",x"AF",x"32",x"20",x"EC",x"32",x"21", -- 0x2E60
		x"EC",x"32",x"22",x"EC",x"CD",x"A7",x"02",x"CD", -- 0x2E68
		x"E0",x"11",x"21",x"00",x"00",x"22",x"02",x"C8", -- 0x2E70
		x"CD",x"16",x"AF",x"CD",x"03",x"AF",x"21",x"9F", -- 0x2E78
		x"B8",x"CD",x"22",x"02",x"CD",x"11",x"B7",x"CD", -- 0x2E80
		x"75",x"B7",x"CD",x"21",x"AF",x"3A",x"01",x"C0", -- 0x2E88
		x"2F",x"32",x"23",x"EC",x"E6",x"10",x"28",x"20", -- 0x2E90
		x"CD",x"16",x"AF",x"CD",x"03",x"AF",x"3A",x"20", -- 0x2E98
		x"EC",x"CD",x"F7",x"66",x"41",x"AF",x"87",x"B5", -- 0x2EA0
		x"7E",x"B3",x"3C",x"B4",x"C7",x"B4",x"59",x"B5", -- 0x2EA8
		x"A3",x"AF",x"DB",x"AF",x"76",x"B0",x"7E",x"B2", -- 0x2EB0
		x"3A",x"22",x"EC",x"B7",x"28",x"03",x"3D",x"18", -- 0x2EB8
		x"3A",x"3A",x"20",x"EC",x"67",x"3A",x"23",x"EC", -- 0x2EC0
		x"E6",x"0C",x"28",x"32",x"E6",x"04",x"20",x"0C", -- 0x2EC8
		x"7C",x"B7",x"28",x"04",x"6C",x"2D",x"18",x"0F", -- 0x2ED0
		x"2E",x"09",x"18",x"0B",x"7C",x"FE",x"09",x"38", -- 0x2ED8
		x"04",x"AF",x"6F",x"18",x"02",x"6C",x"2C",x"22", -- 0x2EE0
		x"20",x"EC",x"CD",x"21",x"AF",x"CD",x"11",x"B7", -- 0x2EE8
		x"CD",x"75",x"B7",x"3A",x"20",x"EC",x"32",x"21", -- 0x2EF0
		x"EC",x"3E",x"06",x"32",x"22",x"EC",x"06",x"02", -- 0x2EF8
		x"DF",x"18",x"8A",x"21",x"40",x"D0",x"16",x"30", -- 0x2F00
		x"CD",x"10",x"AF",x"16",x"00",x"21",x"40",x"D4", -- 0x2F08
		x"01",x"20",x"1C",x"C3",x"53",x"02",x"06",x"02", -- 0x2F10
		x"DF",x"3A",x"01",x"C0",x"E6",x"10",x"28",x"F6", -- 0x2F18
		x"C9",x"2A",x"20",x"EC",x"0E",x"00",x"CD",x"2C", -- 0x2F20
		x"AF",x"65",x"0E",x"16",x"E5",x"11",x"60",x"D4", -- 0x2F28
		x"3E",x"1A",x"CB",x"04",x"94",x"6F",x"26",x"00", -- 0x2F30
		x"19",x"71",x"11",x"20",x"00",x"19",x"71",x"E1", -- 0x2F38
		x"C9",x"21",x"49",x"B9",x"CD",x"22",x"02",x"21", -- 0x2F40
		x"18",x"D1",x"11",x"32",x"B8",x"01",x"05",x"07", -- 0x2F48
		x"CD",x"17",x"AE",x"21",x"78",x"D1",x"01",x"00", -- 0x2F50
		x"05",x"CD",x"34",x"AE",x"CD",x"4B",x"B7",x"CD", -- 0x2F58
		x"75",x"B7",x"3A",x"01",x"C0",x"2F",x"E6",x"1F", -- 0x2F60
		x"FE",x"11",x"30",x"1A",x"DD",x"21",x"18",x"D2", -- 0x2F68
		x"FD",x"21",x"00",x"C0",x"06",x"05",x"CD",x"8C", -- 0x2F70
		x"AF",x"FD",x"23",x"DD",x"2B",x"DD",x"2B",x"10", -- 0x2F78
		x"F5",x"06",x"03",x"DF",x"18",x"DC",x"06",x"14", -- 0x2F80
		x"DF",x"C3",x"6C",x"AE",x"FD",x"7E",x"00",x"DD", -- 0x2F88
		x"E5",x"E1",x"0E",x"08",x"07",x"16",x"00",x"38", -- 0x2F90
		x"01",x"14",x"72",x"11",x"20",x"00",x"19",x"0D", -- 0x2F98
		x"20",x"F2",x"C9",x"21",x"6A",x"B9",x"CD",x"22", -- 0x2FA0
		x"02",x"CD",x"2B",x"B7",x"CD",x"75",x"B7",x"21", -- 0x2FA8
		x"21",x"D1",x"CD",x"79",x"B7",x"21",x"40",x"D5", -- 0x2FB0
		x"01",x"00",x"01",x"16",x"3E",x"CD",x"E2",x"01", -- 0x2FB8
		x"01",x"00",x"01",x"16",x"BE",x"CD",x"E2",x"01", -- 0x2FC0
		x"21",x"40",x"D1",x"CD",x"D4",x"AF",x"CD",x"D4", -- 0x2FC8
		x"AF",x"C3",x"7A",x"B5",x"AF",x"77",x"23",x"3C", -- 0x2FD0
		x"20",x"FB",x"C9",x"21",x"B3",x"B9",x"CD",x"22", -- 0x2FD8
		x"02",x"CD",x"58",x"B7",x"CD",x"75",x"B7",x"AF", -- 0x2FE0
		x"32",x"30",x"EC",x"CD",x"17",x"B0",x"06",x"02", -- 0x2FE8
		x"DF",x"3A",x"01",x"C0",x"2F",x"4F",x"E6",x"10", -- 0x2FF0
		x"C2",x"86",x"AF",x"79",x"E6",x"03",x"28",x"EE", -- 0x2FF8
		x"21",x"30",x"EC",x"E6",x"02",x"3E",x"FF",x"20", -- 0x3000
		x"02",x"3E",x"01",x"86",x"E6",x"07",x"77",x"CD", -- 0x3008
		x"17",x"B0",x"06",x"08",x"DF",x"18",x"D7",x"3A", -- 0x3010
		x"30",x"EC",x"E6",x"07",x"0F",x"0F",x"5F",x"E6", -- 0x3018
		x"01",x"57",x"CB",x"83",x"D5",x"21",x"64",x"D0", -- 0x3020
		x"06",x"04",x"C5",x"CD",x"66",x"B0",x"23",x"23", -- 0x3028
		x"CD",x"66",x"B0",x"23",x"23",x"23",x"23",x"C1", -- 0x3030
		x"10",x"F0",x"D1",x"CB",x"0A",x"21",x"45",x"D8", -- 0x3038
		x"06",x"04",x"C5",x"CD",x"50",x"B0",x"CD",x"50", -- 0x3040
		x"B0",x"0E",x"20",x"09",x"C1",x"10",x"F3",x"C9", -- 0x3048
		x"06",x"08",x"73",x"CB",x"E5",x"7A",x"E6",x"80", -- 0x3050
		x"F6",x"1E",x"77",x"CB",x"A5",x"23",x"13",x"10", -- 0x3058
		x"F1",x"01",x"18",x"00",x"09",x"C9",x"E5",x"7A", -- 0x3060
		x"CD",x"0F",x"AE",x"7B",x"CD",x"06",x"AE",x"21", -- 0x3068
		x"08",x"00",x"19",x"EB",x"E1",x"C9",x"21",x"C1", -- 0x3070
		x"B9",x"CD",x"22",x"02",x"AF",x"32",x"30",x"EC", -- 0x3078
		x"21",x"56",x"B2",x"11",x"40",x"EC",x"CD",x"25", -- 0x3080
		x"B2",x"21",x"57",x"B2",x"11",x"50",x"EC",x"CD", -- 0x3088
		x"35",x"B2",x"21",x"79",x"D0",x"CD",x"6F",x"B1", -- 0x3090
		x"2B",x"2B",x"CD",x"6F",x"B1",x"2B",x"2B",x"CD", -- 0x3098
		x"6F",x"B1",x"CD",x"6F",x"B1",x"2B",x"2B",x"CD", -- 0x30A0
		x"6F",x"B1",x"CD",x"6F",x"B1",x"CD",x"E2",x"B1", -- 0x30A8
		x"CD",x"58",x"B7",x"CD",x"75",x"B7",x"21",x"56", -- 0x30B0
		x"B2",x"11",x"00",x"EB",x"01",x"28",x"00",x"ED", -- 0x30B8
		x"B0",x"CD",x"55",x"B1",x"CD",x"80",x"B1",x"3A", -- 0x30C0
		x"01",x"C0",x"2F",x"4F",x"E6",x"10",x"C2",x"86", -- 0x30C8
		x"AF",x"79",x"E6",x"0F",x"28",x"79",x"E6",x"0C", -- 0x30D0
		x"28",x"2A",x"E6",x"08",x"28",x"16",x"CD",x"59", -- 0x30D8
		x"B1",x"21",x"30",x"EC",x"7E",x"B7",x"20",x"02", -- 0x30E0
		x"3E",x"0C",x"3D",x"77",x"CD",x"55",x"B1",x"06", -- 0x30E8
		x"08",x"DF",x"18",x"58",x"CD",x"59",x"B1",x"21", -- 0x30F0
		x"30",x"EC",x"7E",x"FE",x"0B",x"38",x"02",x"3E", -- 0x30F8
		x"FF",x"3C",x"18",x"E7",x"06",x"FF",x"21",x"40", -- 0x3100
		x"EC",x"3A",x"30",x"EC",x"0F",x"30",x"05",x"06", -- 0x3108
		x"0F",x"21",x"50",x"EC",x"E6",x"07",x"5F",x"16", -- 0x3110
		x"00",x"19",x"79",x"0E",x"00",x"E6",x"02",x"7E", -- 0x3118
		x"57",x"28",x"08",x"3D",x"FE",x"FF",x"20",x"08", -- 0x3120
		x"0C",x"18",x"05",x"3C",x"B7",x"20",x"01",x"0C", -- 0x3128
		x"A0",x"77",x"78",x"3C",x"20",x"0E",x"79",x"B7", -- 0x3130
		x"28",x"0F",x"CB",x"E5",x"7E",x"EE",x"20",x"77", -- 0x3138
		x"CB",x"A5",x"18",x"05",x"7A",x"E6",x"20",x"B6", -- 0x3140
		x"77",x"CD",x"80",x"B1",x"06",x"0A",x"DF",x"06", -- 0x3148
		x"02",x"DF",x"C3",x"C7",x"B0",x"0E",x"16",x"18", -- 0x3150
		x"02",x"0E",x"00",x"21",x"B0",x"B7",x"3A",x"30", -- 0x3158
		x"EC",x"07",x"5F",x"16",x"00",x"19",x"5E",x"23", -- 0x3160
		x"56",x"EB",x"06",x"05",x"C3",x"49",x"02",x"11", -- 0x3168
		x"20",x"00",x"36",x"19",x"CD",x"79",x"B1",x"36", -- 0x3170
		x"0C",x"E5",x"19",x"36",x"25",x"E1",x"2B",x"C9", -- 0x3178
		x"CD",x"E2",x"B1",x"DD",x"21",x"40",x"EC",x"21", -- 0x3180
		x"00",x"EB",x"11",x"04",x"00",x"06",x"04",x"CD", -- 0x3188
		x"C6",x"B1",x"06",x"02",x"CD",x"C6",x"B1",x"06", -- 0x3190
		x"04",x"DD",x"7E",x"00",x"77",x"19",x"DD",x"23", -- 0x3198
		x"10",x"F7",x"DD",x"21",x"50",x"EC",x"21",x"01", -- 0x31A0
		x"EB",x"06",x"04",x"CD",x"D1",x"B1",x"06",x"02", -- 0x31A8
		x"CD",x"D1",x"B1",x"06",x"04",x"DD",x"7E",x"00", -- 0x31B0
		x"E6",x"2F",x"4F",x"7E",x"E6",x"C0",x"B1",x"77", -- 0x31B8
		x"19",x"DD",x"23",x"10",x"F0",x"C9",x"DD",x"7E", -- 0x31C0
		x"00",x"77",x"3C",x"19",x"10",x"FB",x"DD",x"23", -- 0x31C8
		x"C9",x"DD",x"7E",x"00",x"E6",x"2F",x"4F",x"7E", -- 0x31D0
		x"E6",x"C0",x"B1",x"77",x"19",x"10",x"F8",x"DD", -- 0x31D8
		x"23",x"C9",x"11",x"40",x"EC",x"21",x"B9",x"D0", -- 0x31E0
		x"CD",x"FD",x"B1",x"2B",x"2B",x"CD",x"FD",x"B1", -- 0x31E8
		x"2B",x"2B",x"CD",x"FD",x"B1",x"CD",x"FD",x"B1", -- 0x31F0
		x"2B",x"2B",x"CD",x"FD",x"B1",x"CB",x"E3",x"1A", -- 0x31F8
		x"CB",x"A3",x"E6",x"20",x"28",x"02",x"3E",x"01", -- 0x3200
		x"CD",x"0F",x"AE",x"CD",x"1C",x"B2",x"CB",x"E3", -- 0x3208
		x"1A",x"CD",x"0F",x"AE",x"CB",x"A3",x"01",x"9F", -- 0x3210
		x"FF",x"09",x"13",x"C9",x"1A",x"CD",x"06",x"AE", -- 0x3218
		x"01",x"DF",x"FF",x"09",x"C9",x"ED",x"A0",x"01", -- 0x3220
		x"0F",x"00",x"09",x"ED",x"A0",x"01",x"07",x"00", -- 0x3228
		x"09",x"0E",x"FF",x"18",x"14",x"7E",x"E6",x"0F", -- 0x3230
		x"12",x"13",x"01",x"10",x"00",x"09",x"7E",x"E6", -- 0x3238
		x"0F",x"12",x"13",x"01",x"08",x"00",x"09",x"0E", -- 0x3240
		x"0F",x"06",x"04",x"7E",x"A1",x"12",x"23",x"23", -- 0x3248
		x"23",x"23",x"13",x"10",x"F6",x"C9",x"00",x"00", -- 0x3250
		x"80",x"C0",x"01",x"00",x"98",x"C0",x"02",x"00", -- 0x3258
		x"B0",x"C0",x"03",x"00",x"C8",x"C0",x"B0",x"40", -- 0x3260
		x"80",x"A0",x"B2",x"40",x"B0",x"A0",x"E0",x"40", -- 0x3268
		x"80",x"80",x"E8",x"40",x"80",x"70",x"80",x"80", -- 0x3270
		x"80",x"50",x"84",x"40",x"90",x"40",x"21",x"50", -- 0x3278
		x"BA",x"CD",x"22",x"02",x"CD",x"65",x"B7",x"CD", -- 0x3280
		x"75",x"B7",x"CD",x"FD",x"2C",x"3E",x"80",x"32", -- 0x3288
		x"00",x"E0",x"CD",x"6A",x"B3",x"21",x"00",x"00", -- 0x3290
		x"22",x"60",x"EC",x"22",x"62",x"EC",x"CD",x"3D", -- 0x3298
		x"B3",x"3A",x"01",x"C0",x"57",x"2F",x"E6",x"1F", -- 0x32A0
		x"FE",x"11",x"D2",x"52",x"B3",x"7A",x"CB",x"67", -- 0x32A8
		x"CA",x"21",x"B3",x"3E",x"00",x"32",x"61",x"EC", -- 0x32B0
		x"7A",x"CB",x"47",x"CA",x"F9",x"B2",x"3E",x"00", -- 0x32B8
		x"32",x"62",x"EC",x"7A",x"CB",x"4F",x"C2",x"F1", -- 0x32C0
		x"B2",x"3A",x"63",x"EC",x"3C",x"32",x"63",x"EC", -- 0x32C8
		x"FE",x"01",x"CA",x"DF",x"B2",x"FE",x"0A",x"C2", -- 0x32D0
		x"37",x"B3",x"3E",x"01",x"32",x"63",x"EC",x"CD", -- 0x32D8
		x"6A",x"B3",x"3A",x"60",x"EC",x"3D",x"E6",x"1F", -- 0x32E0
		x"32",x"60",x"EC",x"CD",x"3D",x"B3",x"C3",x"37", -- 0x32E8
		x"B3",x"3E",x"00",x"32",x"63",x"EC",x"C3",x"37", -- 0x32F0
		x"B3",x"3A",x"62",x"EC",x"3C",x"32",x"62",x"EC", -- 0x32F8
		x"FE",x"01",x"CA",x"0F",x"B3",x"FE",x"0A",x"C2", -- 0x3300
		x"37",x"B3",x"3E",x"01",x"32",x"62",x"EC",x"CD", -- 0x3308
		x"6A",x"B3",x"3A",x"60",x"EC",x"3C",x"E6",x"1F", -- 0x3310
		x"32",x"60",x"EC",x"CD",x"3D",x"B3",x"C3",x"37", -- 0x3318
		x"B3",x"3A",x"61",x"EC",x"FE",x"00",x"C2",x"37", -- 0x3320
		x"B3",x"3A",x"60",x"EC",x"4F",x"CD",x"78",x"11", -- 0x3328
		x"3A",x"61",x"EC",x"3C",x"32",x"61",x"EC",x"06", -- 0x3330
		x"02",x"DF",x"C3",x"A1",x"B2",x"3A",x"60",x"EC", -- 0x3338
		x"E6",x"0F",x"32",x"D0",x"D2",x"3A",x"60",x"EC", -- 0x3340
		x"07",x"07",x"07",x"07",x"E6",x"0F",x"32",x"B0", -- 0x3348
		x"D2",x"C9",x"CD",x"6A",x"B3",x"CD",x"FD",x"2C", -- 0x3350
		x"AF",x"32",x"00",x"E0",x"06",x"02",x"DF",x"3A", -- 0x3358
		x"01",x"C0",x"2F",x"E6",x"1F",x"20",x"F5",x"C3", -- 0x3360
		x"86",x"AF",x"0E",x"00",x"CD",x"78",x"11",x"0E", -- 0x3368
		x"0B",x"CD",x"78",x"11",x"0E",x"10",x"CD",x"78", -- 0x3370
		x"11",x"0E",x"0F",x"C3",x"78",x"11",x"CD",x"2B", -- 0x3378
		x"B7",x"CD",x"75",x"B7",x"21",x"22",x"BA",x"CD", -- 0x3380
		x"22",x"02",x"21",x"68",x"D0",x"CD",x"31",x"B4", -- 0x3388
		x"21",x"E8",x"D0",x"CD",x"33",x"B4",x"21",x"68", -- 0x3390
		x"D1",x"CD",x"31",x"B4",x"21",x"28",x"D2",x"CD", -- 0x3398
		x"33",x"B4",x"21",x"E5",x"D2",x"01",x"00",x"04", -- 0x33A0
		x"CD",x"24",x"B4",x"CD",x"24",x"B4",x"23",x"10", -- 0x33A8
		x"F7",x"DD",x"21",x"C8",x"B7",x"FD",x"21",x"88", -- 0x33B0
		x"D0",x"CD",x"E1",x"B3",x"FD",x"21",x"08",x"D1", -- 0x33B8
		x"CD",x"E1",x"B3",x"DD",x"21",x"E8",x"B7",x"21", -- 0x33C0
		x"86",x"D8",x"CD",x"07",x"B4",x"21",x"89",x"D8", -- 0x33C8
		x"CD",x"07",x"B4",x"21",x"08",x"B8",x"11",x"00", -- 0x33D0
		x"EB",x"01",x"20",x"00",x"ED",x"B0",x"C3",x"7A", -- 0x33D8
		x"B5",x"06",x"08",x"C5",x"CD",x"F9",x"B3",x"FD", -- 0x33E0
		x"E5",x"E1",x"01",x"00",x"04",x"09",x"CD",x"FC", -- 0x33E8
		x"B3",x"C1",x"FD",x"23",x"FD",x"23",x"10",x"EB", -- 0x33F0
		x"C9",x"FD",x"E5",x"E1",x"01",x"02",x"02",x"DD", -- 0x33F8
		x"56",x"00",x"DD",x"23",x"C3",x"53",x"02",x"06", -- 0x3400
		x"08",x"C5",x"CD",x"1A",x"B4",x"CB",x"E5",x"CD", -- 0x3408
		x"1A",x"B4",x"01",x"10",x"00",x"09",x"C1",x"10", -- 0x3410
		x"F0",x"C9",x"DD",x"56",x"00",x"72",x"23",x"72", -- 0x3418
		x"2B",x"DD",x"23",x"C9",x"71",x"0C",x"11",x"C0", -- 0x3420
		x"00",x"19",x"71",x"0C",x"11",x"42",x"FF",x"19", -- 0x3428
		x"C9",x"0E",x"00",x"06",x"08",x"71",x"0C",x"23", -- 0x3430
		x"23",x"10",x"FA",x"C9",x"21",x"A8",x"BA",x"CD", -- 0x3438
		x"22",x"02",x"CD",x"2B",x"B7",x"CD",x"75",x"B7", -- 0x3440
		x"21",x"B7",x"D0",x"06",x"0F",x"70",x"2B",x"10", -- 0x3448
		x"FC",x"70",x"21",x"F9",x"D0",x"11",x"20",x"00", -- 0x3450
		x"06",x"04",x"36",x"50",x"19",x"36",x"53",x"19", -- 0x3458
		x"36",x"54",x"19",x"36",x"57",x"19",x"19",x"10", -- 0x3460
		x"F1",x"21",x"E8",x"D0",x"CD",x"9E",x"B4",x"21", -- 0x3468
		x"88",x"D1",x"CD",x"9E",x"B4",x"21",x"28",x"D2", -- 0x3470
		x"CD",x"9E",x"B4",x"21",x"C8",x"D2",x"CD",x"9E", -- 0x3478
		x"B4",x"0E",x"00",x"21",x"E8",x"D4",x"CD",x"B4", -- 0x3480
		x"B4",x"21",x"88",x"D5",x"CD",x"B4",x"B4",x"21", -- 0x3488
		x"28",x"D6",x"CD",x"B4",x"B4",x"21",x"C8",x"D6", -- 0x3490
		x"CD",x"B4",x"B4",x"C3",x"7A",x"B5",x"06",x"10", -- 0x3498
		x"C5",x"E5",x"3E",x"30",x"06",x"04",x"11",x"20", -- 0x34A0
		x"00",x"77",x"19",x"3C",x"10",x"FB",x"E1",x"23", -- 0x34A8
		x"C1",x"10",x"ED",x"C9",x"06",x"10",x"E5",x"3E", -- 0x34B0
		x"04",x"71",x"11",x"20",x"00",x"19",x"3D",x"20", -- 0x34B8
		x"F8",x"E1",x"0C",x"23",x"10",x"F0",x"C9",x"CD", -- 0x34C0
		x"58",x"B7",x"CD",x"75",x"B7",x"21",x"C1",x"BA", -- 0x34C8
		x"CD",x"22",x"02",x"AF",x"32",x"30",x"EC",x"21", -- 0x34D0
		x"85",x"D8",x"0E",x"F8",x"CD",x"40",x"B5",x"CD", -- 0x34D8
		x"0B",x"B5",x"06",x"02",x"DF",x"3A",x"01",x"C0", -- 0x34E0
		x"2F",x"4F",x"E6",x"10",x"C2",x"86",x"AF",x"79", -- 0x34E8
		x"E6",x"03",x"28",x"EE",x"21",x"30",x"EC",x"E6", -- 0x34F0
		x"02",x"3E",x"FF",x"20",x"02",x"3E",x"01",x"86", -- 0x34F8
		x"E6",x"03",x"77",x"CD",x"0B",x"B5",x"06",x"08", -- 0x3500
		x"DF",x"18",x"D7",x"21",x"88",x"D0",x"3A",x"30", -- 0x3508
		x"EC",x"E6",x"02",x"0F",x"4F",x"06",x"08",x"71", -- 0x3510
		x"23",x"23",x"10",x"FB",x"21",x"A8",x"D0",x"3A", -- 0x3518
		x"30",x"EC",x"E6",x"01",x"28",x"02",x"3E",x"08", -- 0x3520
		x"4F",x"06",x"08",x"71",x"23",x"23",x"0C",x"10", -- 0x3528
		x"FA",x"3A",x"30",x"EC",x"E6",x"03",x"07",x"07", -- 0x3530
		x"07",x"F6",x"80",x"4F",x"3C",x"21",x"95",x"D8", -- 0x3538
		x"06",x"08",x"C5",x"E5",x"71",x"23",x"B7",x"20", -- 0x3540
		x"01",x"0C",x"10",x"F8",x"E1",x"01",x"20",x"00", -- 0x3548
		x"09",x"C1",x"B7",x"28",x"01",x"0C",x"10",x"EA", -- 0x3550
		x"C9",x"16",x"3C",x"CD",x"0D",x"AF",x"0E",x"0E", -- 0x3558
		x"21",x"40",x"D0",x"06",x"10",x"36",x"4C",x"23", -- 0x3560
		x"36",x"4D",x"23",x"10",x"F8",x"06",x"10",x"36", -- 0x3568
		x"4E",x"23",x"36",x"4F",x"23",x"10",x"F8",x"0D", -- 0x3570
		x"20",x"E9",x"06",x"02",x"DF",x"3A",x"01",x"C0", -- 0x3578
		x"E6",x"10",x"20",x"F6",x"C3",x"86",x"AF",x"21", -- 0x3580
		x"6F",x"BA",x"CD",x"22",x"02",x"21",x"18",x"D1", -- 0x3588
		x"11",x"39",x"B8",x"01",x"07",x"07",x"CD",x"17", -- 0x3590
		x"AE",x"21",x"78",x"D1",x"01",x"00",x"07",x"CD", -- 0x3598
		x"34",x"AE",x"CD",x"3B",x"B7",x"CD",x"75",x"B7", -- 0x35A0
		x"AF",x"67",x"6F",x"22",x"2A",x"EC",x"22",x"2C", -- 0x35A8
		x"EC",x"32",x"22",x"EC",x"32",x"2E",x"EC",x"21", -- 0x35B0
		x"34",x"EC",x"CD",x"B2",x"AD",x"2B",x"36",x"02", -- 0x35B8
		x"21",x"2C",x"EC",x"06",x"07",x"C5",x"E5",x"CD", -- 0x35C0
		x"AA",x"B6",x"E1",x"34",x"C1",x"10",x"F6",x"70", -- 0x35C8
		x"CD",x"E0",x"B6",x"3A",x"01",x"C0",x"2F",x"4F", -- 0x35D0
		x"E6",x"1F",x"FE",x"11",x"D2",x"94",x"B6",x"3A", -- 0x35D8
		x"24",x"EC",x"B7",x"28",x"03",x"3D",x"18",x"46", -- 0x35E0
		x"3A",x"2E",x"EC",x"B7",x"79",x"20",x"0F",x"E6", -- 0x35E8
		x"10",x"28",x"40",x"AF",x"32",x"2F",x"EC",x"3C", -- 0x35F0
		x"32",x"2E",x"EC",x"C3",x"8E",x"B6",x"E6",x"10", -- 0x35F8
		x"20",x"31",x"32",x"2E",x"EC",x"0E",x"80",x"3A", -- 0x3600
		x"2A",x"EC",x"B7",x"28",x"05",x"CB",x"09",x"3D", -- 0x3608
		x"18",x"F8",x"21",x"34",x"EC",x"3A",x"2C",x"EC", -- 0x3610
		x"5F",x"16",x"00",x"19",x"FE",x"06",x"7E",x"20", -- 0x3618
		x"06",x"79",x"E6",x"03",x"7E",x"20",x"02",x"A9", -- 0x3620
		x"77",x"CD",x"AA",x"B6",x"3E",x"03",x"32",x"24", -- 0x3628
		x"EC",x"18",x"5B",x"3A",x"22",x"EC",x"B7",x"28", -- 0x3630
		x"03",x"3D",x"18",x"4F",x"79",x"E6",x"03",x"28", -- 0x3638
		x"1B",x"E6",x"02",x"3A",x"2A",x"EC",x"28",x"08", -- 0x3640
		x"B7",x"20",x"02",x"3E",x"08",x"3D",x"18",x"07", -- 0x3648
		x"FE",x"07",x"38",x"02",x"3E",x"FF",x"3C",x"32", -- 0x3650
		x"2A",x"EC",x"18",x"1E",x"79",x"E6",x"0C",x"28", -- 0x3658
		x"2D",x"E6",x"08",x"3A",x"2C",x"EC",x"28",x"08", -- 0x3660
		x"B7",x"20",x"02",x"3E",x"07",x"3D",x"18",x"07", -- 0x3668
		x"FE",x"06",x"38",x"02",x"3E",x"FF",x"3C",x"32", -- 0x3670
		x"2C",x"EC",x"CD",x"E0",x"B6",x"3A",x"2A",x"EC", -- 0x3678
		x"32",x"2B",x"EC",x"3A",x"2C",x"EC",x"32",x"2D", -- 0x3680
		x"EC",x"3E",x"03",x"32",x"22",x"EC",x"06",x"02", -- 0x3688
		x"DF",x"C3",x"D3",x"B5",x"AF",x"32",x"22",x"EC", -- 0x3690
		x"32",x"24",x"EC",x"21",x"34",x"EC",x"CD",x"B2", -- 0x3698
		x"AD",x"2B",x"36",x"02",x"CD",x"AA",x"B6",x"C3", -- 0x36A0
		x"86",x"AF",x"21",x"34",x"EC",x"3A",x"2C",x"EC", -- 0x36A8
		x"5F",x"16",x"00",x"19",x"FE",x"06",x"7E",x"20", -- 0x36B0
		x"04",x"E6",x"FC",x"F6",x"02",x"4F",x"CD",x"04", -- 0x36B8
		x"B7",x"11",x"00",x"FC",x"19",x"11",x"20",x"00", -- 0x36C0
		x"06",x"08",x"AF",x"CB",x"01",x"30",x"01",x"3C", -- 0x36C8
		x"77",x"19",x"10",x"F6",x"21",x"34",x"EC",x"11", -- 0x36D0
		x"00",x"C8",x"01",x"07",x"00",x"ED",x"B0",x"C9", -- 0x36D8
		x"3A",x"2B",x"EC",x"47",x"3A",x"2D",x"EC",x"0E", -- 0x36E0
		x"00",x"CD",x"F5",x"B6",x"3A",x"2A",x"EC",x"47", -- 0x36E8
		x"3A",x"2C",x"EC",x"0E",x"16",x"CD",x"07",x"B7", -- 0x36F0
		x"EB",x"68",x"26",x"00",x"29",x"29",x"29",x"29", -- 0x36F8
		x"29",x"19",x"71",x"C9",x"3A",x"2C",x"EC",x"21", -- 0x3700
		x"18",x"D6",x"B7",x"C8",x"2B",x"2B",x"3D",x"18", -- 0x3708
		x"FA",x"06",x"06",x"11",x"F5",x"BA",x"21",x"60", -- 0x3710
		x"D0",x"C3",x"EE",x"01",x"11",x"05",x"BB",x"06", -- 0x3718
		x"01",x"C3",x"EE",x"01",x"11",x"FB",x"BA",x"06", -- 0x3720
		x"0A",x"18",x"EB",x"21",x"60",x"D0",x"11",x"06", -- 0x3728
		x"BB",x"06",x"05",x"C3",x"EE",x"01",x"CD",x"1C", -- 0x3730
		x"B7",x"18",x"F3",x"21",x"60",x"D0",x"06",x"08", -- 0x3738
		x"11",x"0B",x"BB",x"CD",x"EE",x"01",x"CD",x"1C", -- 0x3740
		x"B7",x"18",x"03",x"21",x"60",x"D0",x"06",x"06", -- 0x3748
		x"11",x"13",x"BB",x"CD",x"EE",x"01",x"18",x"D6", -- 0x3750
		x"21",x"60",x"D0",x"06",x"0D",x"11",x"19",x"BB", -- 0x3758
		x"CD",x"EE",x"01",x"18",x"D1",x"21",x"60",x"D0", -- 0x3760
		x"06",x"0D",x"11",x"19",x"BB",x"CD",x"EE",x"01", -- 0x3768
		x"CD",x"1C",x"B7",x"18",x"D9",x"01",x"85",x"B7", -- 0x3770
		x"C5",x"01",x"20",x"00",x"7C",x"FE",x"D4",x"D0", -- 0x3778
		x"36",x"30",x"09",x"18",x"F7",x"21",x"41",x"D0", -- 0x3780
		x"16",x"35",x"01",x"01",x"1C",x"C3",x"53",x"02", -- 0x3788
		x"60",x"80",x"C0",x"00",x"C0",x"00",x"40",x"80", -- 0x3790
		x"00",x"01",x"20",x"01",x"50",x"00",x"60",x"80", -- 0x3798
		x"20",x"80",x"30",x"00",x"38",x"80",x"30",x"00", -- 0x37A0
		x"30",x"00",x"38",x"00",x"28",x"00",x"60",x"80", -- 0x37A8
		x"79",x"D4",x"78",x"D4",x"75",x"D4",x"74",x"D4", -- 0x37B0
		x"71",x"D4",x"70",x"D4",x"6F",x"D4",x"6E",x"D4", -- 0x37B8
		x"6B",x"D4",x"6A",x"D4",x"69",x"D4",x"68",x"D4", -- 0x37C0
		x"31",x"10",x"31",x"11",x"31",x"12",x"31",x"13", -- 0x37C8
		x"31",x"14",x"31",x"15",x"31",x"16",x"31",x"17", -- 0x37D0
		x"31",x"18",x"31",x"19",x"31",x"1A",x"31",x"1B", -- 0x37D8
		x"31",x"1C",x"31",x"1D",x"31",x"1E",x"31",x"1F", -- 0x37E0
		x"F8",x"9E",x"F9",x"9E",x"FA",x"9E",x"FB",x"9E", -- 0x37E8
		x"FC",x"9E",x"FD",x"9E",x"FE",x"9E",x"FF",x"9E", -- 0x37F0
		x"FA",x"9F",x"FB",x"9F",x"FC",x"9F",x"FD",x"9F", -- 0x37F8
		x"FE",x"9F",x"F9",x"9F",x"FF",x"9F",x"FF",x"90", -- 0x3800
		x"70",x"66",x"C4",x"28",x"72",x"66",x"C4",x"38", -- 0x3808
		x"74",x"66",x"C4",x"50",x"76",x"66",x"C4",x"60", -- 0x3810
		x"78",x"66",x"C4",x"78",x"7A",x"66",x"C4",x"88", -- 0x3818
		x"7C",x"66",x"C4",x"A0",x"7E",x"66",x"C4",x"B0", -- 0x3820
		x"25",x"18",x"14",x"25",x"30",x"4B",x"4B",x"30", -- 0x3828
		x"4B",x"4B",x"0C",x"00",x"00",x"00",x"11",x"30", -- 0x3830
		x"44",x"0C",x"08",x"00",x"00",x"11",x"30",x"44", -- 0x3838
		x"03",x"17",x"00",x"09",x"03",x"17",x"01",x"00", -- 0x3840
		x"03",x"0D",x"00",x"02",x"03",x"0A",x"00",x"09", -- 0x3848
		x"00",x"0D",x"3C",x"D1",x"48",x"30",x"1B",x"0A", -- 0x3850
		x"16",x"30",x"0C",x"11",x"0E",x"0C",x"14",x"30", -- 0x3858
		x"49",x"0F",x"B6",x"D1",x"0A",x"0D",x"0D",x"1B", -- 0x3860
		x"30",x"20",x"1B",x"30",x"1B",x"0D",x"30",x"30", -- 0x3868
		x"15",x"18",x"0C",x"08",x"94",x"D0",x"20",x"25", -- 0x3870
		x"1B",x"0A",x"16",x"01",x"30",x"44",x"08",x"92", -- 0x3878
		x"D0",x"20",x"25",x"1B",x"0A",x"16",x"02",x"30", -- 0x3880
		x"44",x"08",x"90",x"D0",x"1F",x"25",x"1B",x"0A", -- 0x3888
		x"16",x"30",x"30",x"44",x"08",x"8E",x"D0",x"1C", -- 0x3890
		x"25",x"1B",x"0A",x"16",x"30",x"30",x"44",x"00", -- 0x3898
		x"0D",x"5E",x"D1",x"48",x"30",x"1D",x"0E",x"1C", -- 0x38A0
		x"1D",x"30",x"16",x"0E",x"17",x"1E",x"30",x"49", -- 0x38A8
		x"08",x"7A",x"D0",x"00",x"01",x"30",x"12",x"17", -- 0x38B0
		x"19",x"1E",x"1D",x"09",x"78",x"D0",x"00",x"02", -- 0x38B8
		x"30",x"18",x"1E",x"1D",x"19",x"1E",x"1D",x"0D", -- 0x38C0
		x"76",x"D0",x"00",x"03",x"30",x"11",x"0A",x"1B", -- 0x38C8
		x"0D",x"30",x"0C",x"18",x"15",x"18",x"1B",x"14", -- 0x38D0
		x"74",x"D0",x"00",x"04",x"30",x"1C",x"18",x"0F", -- 0x38D8
		x"1D",x"30",x"0C",x"18",x"15",x"18",x"1B",x"30", -- 0x38E0
		x"44",x"30",x"0C",x"11",x"0A",x"1B",x"16",x"72", -- 0x38E8
		x"D0",x"00",x"05",x"30",x"1C",x"18",x"0F",x"1D", -- 0x38F0
		x"30",x"0C",x"18",x"15",x"18",x"1B",x"30",x"44", -- 0x38F8
		x"30",x"1C",x"0C",x"1B",x"18",x"15",x"15",x"12", -- 0x3900
		x"70",x"D0",x"00",x"06",x"30",x"0D",x"18",x"1D", -- 0x3908
		x"30",x"0C",x"1B",x"18",x"1C",x"1C",x"30",x"11", -- 0x3910
		x"0A",x"1D",x"0C",x"11",x"07",x"6E",x"D0",x"00", -- 0x3918
		x"07",x"30",x"0C",x"11",x"0A",x"1B",x"09",x"6C", -- 0x3920
		x"D0",x"00",x"08",x"30",x"1C",x"0C",x"1B",x"18", -- 0x3928
		x"15",x"15",x"09",x"6A",x"D0",x"00",x"09",x"30", -- 0x3930
		x"18",x"0B",x"13",x"0E",x"0C",x"1D",x"08",x"68", -- 0x3938
		x"D0",x"01",x"00",x"30",x"1C",x"18",x"1E",x"17", -- 0x3940
		x"0D",x"00",x"09",x"7D",x"D1",x"48",x"30",x"12", -- 0x3948
		x"17",x"19",x"1E",x"1D",x"30",x"49",x"11",x"FA", -- 0x3950
		x"D0",x"12",x"17",x"25",x"0A",x"0D",x"0D",x"1B", -- 0x3958
		x"30",x"30",x"16",x"1C",x"0B",x"30",x"30",x"15", -- 0x3960
		x"1C",x"0B",x"00",x"02",x"F9",x"D4",x"3E",x"3E", -- 0x3968
		x"02",x"F7",x"D4",x"3E",x"3E",x"02",x"F5",x"D4", -- 0x3970
		x"3E",x"3E",x"02",x"F3",x"D4",x"3E",x"3E",x"02", -- 0x3978
		x"F9",x"D0",x"30",x"30",x"02",x"F7",x"D0",x"31", -- 0x3980
		x"31",x"02",x"F5",x"D0",x"32",x"32",x"02",x"F3", -- 0x3988
		x"D0",x"33",x"33",x"05",x"99",x"D0",x"17",x"18", -- 0x3990
		x"30",x"30",x"30",x"05",x"97",x"D0",x"22",x"30", -- 0x3998
		x"30",x"31",x"31",x"05",x"95",x"D0",x"23",x"30", -- 0x39A0
		x"30",x"32",x"32",x"05",x"93",x"D0",x"22",x"23", -- 0x39A8
		x"30",x"33",x"33",x"00",x"0A",x"7D",x"D1",x"48", -- 0x39B0
		x"30",x"1C",x"0C",x"1B",x"18",x"15",x"15",x"30", -- 0x39B8
		x"49",x"00",x"0A",x"7D",x"D1",x"48",x"30",x"18", -- 0x39C0
		x"0B",x"13",x"0E",x"0C",x"1D",x"30",x"49",x"05", -- 0x39C8
		x"38",x"D1",x"01",x"06",x"21",x"01",x"06",x"05", -- 0x39D0
		x"34",x"D1",x"01",x"06",x"21",x"03",x"02",x"05", -- 0x39D8
		x"30",x"D1",x"01",x"06",x"21",x"03",x"02",x"05", -- 0x39E0
		x"2E",x"D1",x"01",x"06",x"21",x"03",x"02",x"05", -- 0x39E8
		x"2A",x"D1",x"01",x"06",x"21",x"06",x"04",x"05", -- 0x39F0
		x"28",x"D1",x"01",x"06",x"21",x"03",x"02",x"0F", -- 0x39F8
		x"65",x"D0",x"4B",x"30",x"19",x"44",x"19",x"0A", -- 0x3A00
		x"1D",x"1D",x"0E",x"1B",x"17",x"30",x"17",x"18", -- 0x3A08
		x"24",x"0E",x"63",x"D0",x"4B",x"30",x"0C",x"44", -- 0x3A10
		x"0C",x"18",x"15",x"18",x"1B",x"30",x"0C",x"18", -- 0x3A18
		x"0D",x"0E",x"00",x"0E",x"3D",x"D1",x"48",x"30", -- 0x3A20
		x"11",x"0A",x"1B",x"0D",x"30",x"0C",x"18",x"15", -- 0x3A28
		x"18",x"1B",x"30",x"49",x"19",x"99",x"D0",x"25", -- 0x3A30
		x"0C",x"11",x"0A",x"1B",x"25",x"30",x"30",x"25", -- 0x3A38
		x"25",x"1C",x"0C",x"1B",x"18",x"15",x"15",x"25", -- 0x3A40
		x"25",x"30",x"18",x"0B",x"13",x"0E",x"0C",x"1D", -- 0x3A48
		x"00",x"09",x"7D",x"D1",x"48",x"30",x"1C",x"18", -- 0x3A50
		x"1E",x"17",x"0D",x"30",x"49",x"0F",x"30",x"D1", -- 0x3A58
		x"1C",x"18",x"1E",x"17",x"0D",x"30",x"0C",x"18", -- 0x3A60
		x"0D",x"0E",x"30",x"2A",x"00",x"00",x"2B",x"00", -- 0x3A68
		x"0A",x"7D",x"D1",x"48",x"30",x"18",x"1E",x"1D", -- 0x3A70
		x"19",x"1E",x"1D",x"30",x"49",x"12",x"DA",x"D0", -- 0x3A78
		x"18",x"1E",x"1D",x"25",x"0A",x"0D",x"0D",x"1B", -- 0x3A80
		x"30",x"30",x"16",x"1C",x"0B",x"30",x"30",x"15", -- 0x3A88
		x"1C",x"0B",x"13",x"C8",x"D0",x"0C",x"08",x"00", -- 0x3A90
		x"06",x"11",x"30",x"0D",x"01",x"25",x"00",x"30", -- 0x3A98
		x"44",x"30",x"17",x"18",x"30",x"1C",x"0E",x"1D", -- 0x3AA0
		x"00",x"15",x"BD",x"D0",x"48",x"30",x"1C",x"18", -- 0x3AA8
		x"0F",x"1D",x"30",x"0C",x"18",x"15",x"18",x"1B", -- 0x3AB0
		x"30",x"44",x"30",x"0C",x"11",x"0A",x"1B",x"30", -- 0x3AB8
		x"49",x"00",x"17",x"9D",x"D0",x"48",x"30",x"1C", -- 0x3AC0
		x"18",x"0F",x"1D",x"30",x"0C",x"18",x"15",x"18", -- 0x3AC8
		x"1B",x"30",x"44",x"30",x"1C",x"0C",x"1B",x"18", -- 0x3AD0
		x"15",x"15",x"30",x"49",x"15",x"79",x"D0",x"0C", -- 0x3AD8
		x"18",x"0D",x"0E",x"30",x"50",x"30",x"54",x"30", -- 0x3AE0
		x"53",x"30",x"57",x"30",x"52",x"30",x"56",x"30", -- 0x3AE8
		x"59",x"30",x"52",x"57",x"00",x"0F",x"44",x"0E", -- 0x3AF0
		x"21",x"0E",x"0C",x"15",x"0E",x"1F",x"0E",x"1B", -- 0x3AF8
		x"44",x"17",x"0E",x"21",x"1D",x"34",x"0F",x"44", -- 0x3B00
		x"0E",x"17",x"0D",x"0F",x"44",x"18",x"17",x"46", -- 0x3B08
		x"18",x"0F",x"0F",x"15",x"0E",x"1F",x"0E",x"1B", -- 0x3B10
		x"26",x"1B",x"1D",x"44",x"12",x"17",x"0C",x"34", -- 0x3B18
		x"15",x"1D",x"44",x"0D",x"0E",x"0C",x"27",x"C1", -- 0x3B20
		x"FF",x"F7",x"E8",x"92",x"F2",x"91",x"C1",x"A9", -- 0x3B28
		x"20",x"9C",x"45",x"B7",x"EC",x"08",x"A9",x"F2", -- 0x3B30
		x"29",x"AD",x"73",x"5F",x"AD",x"EA",x"FF",x"61", -- 0x3B38
		x"A4",x"02",x"8A",x"80",x"D4",x"18",x"A8",x"DB", -- 0x3B40
		x"A4",x"40",x"46",x"10",x"4F",x"23",x"BA",x"0C", -- 0x3B48
		x"04",x"01",x"AA",x"B3",x"E9",x"B1",x"F3",x"2C", -- 0x3B50
		x"C5",x"D1",x"35",x"82",x"F0",x"00",x"83",x"6C", -- 0x3B58
		x"8A",x"98",x"D2",x"01",x"EB",x"71",x"E6",x"8A", -- 0x3B60
		x"9B",x"90",x"78",x"63",x"36",x"09",x"49",x"10", -- 0x3B68
		x"87",x"23",x"68",x"8D",x"F5",x"73",x"D4",x"C5", -- 0x3B70
		x"E6",x"8F",x"41",x"F0",x"55",x"39",x"69",x"0B", -- 0x3B78
		x"65",x"18",x"31",x"89",x"59",x"A7",x"EF",x"04", -- 0x3B80
		x"9B",x"84",x"E5",x"60",x"33",x"0E",x"6F",x"04", -- 0x3B88
		x"FC",x"7B",x"D4",x"B9",x"7D",x"58",x"7F",x"F6", -- 0x3B90
		x"9E",x"C0",x"6A",x"EA",x"F9",x"30",x"F7",x"0C", -- 0x3B98
		x"A6",x"59",x"D0",x"0A",x"69",x"48",x"E6",x"80", -- 0x3BA0
		x"44",x"48",x"77",x"CD",x"CA",x"AE",x"5F",x"E0", -- 0x3BA8
		x"9A",x"B1",x"EF",x"82",x"9D",x"D8",x"2E",x"E3", -- 0x3BB0
		x"CF",x"57",x"74",x"B0",x"6D",x"3F",x"BA",x"AA", -- 0x3BB8
		x"21",x"40",x"E2",x"11",x"FE",x"01",x"7F",x"68", -- 0x3BC0
		x"B1",x"40",x"84",x"42",x"11",x"24",x"C4",x"85", -- 0x3BC8
		x"F4",x"4C",x"CC",x"48",x"B6",x"2B",x"80",x"8B", -- 0x3BD0
		x"5F",x"C9",x"BF",x"BD",x"F9",x"FA",x"3E",x"99", -- 0x3BD8
		x"99",x"07",x"68",x"90",x"DD",x"EF",x"8C",x"64", -- 0x3BE0
		x"EB",x"A9",x"D6",x"80",x"C7",x"C1",x"00",x"E1", -- 0x3BE8
		x"54",x"0C",x"60",x"C0",x"FB",x"C6",x"67",x"4A", -- 0x3BF0
		x"FF",x"00",x"BA",x"EA",x"AD",x"A6",x"70",x"21", -- 0x3BF8
		x"F4",x"85",x"56",x"88",x"48",x"44",x"BB",x"21", -- 0x3C00
		x"EA",x"48",x"A0",x"13",x"0B",x"21",x"C8",x"12", -- 0x3C08
		x"BE",x"00",x"3D",x"A2",x"DE",x"00",x"45",x"55", -- 0x3C10
		x"26",x"96",x"EF",x"DE",x"19",x"03",x"C8",x"03", -- 0x3C18
		x"D7",x"41",x"1A",x"E1",x"B5",x"85",x"F4",x"22", -- 0x3C20
		x"28",x"69",x"BE",x"63",x"2E",x"77",x"FF",x"D0", -- 0x3C28
		x"45",x"4A",x"9B",x"15",x"CE",x"21",x"F9",x"63", -- 0x3C30
		x"D0",x"9F",x"6A",x"11",x"DD",x"94",x"B2",x"71", -- 0x3C38
		x"B8",x"0B",x"A6",x"91",x"B7",x"44",x"63",x"E2", -- 0x3C40
		x"A0",x"44",x"B3",x"89",x"42",x"41",x"A0",x"88", -- 0x3C48
		x"4B",x"0F",x"60",x"44",x"6F",x"49",x"CD",x"31", -- 0x3C50
		x"39",x"3B",x"BA",x"FA",x"BB",x"F4",x"5A",x"55", -- 0x3C58
		x"96",x"9B",x"B0",x"88",x"32",x"6C",x"26",x"CB", -- 0x3C60
		x"E5",x"E8",x"19",x"0E",x"76",x"C3",x"4E",x"48", -- 0x3C68
		x"1F",x"25",x"D2",x"DF",x"26",x"68",x"EB",x"25", -- 0x3C70
		x"59",x"EA",x"FF",x"50",x"AF",x"93",x"D1",x"93", -- 0x3C78
		x"EF",x"C0",x"0E",x"00",x"E4",x"42",x"3F",x"47", -- 0x3C80
		x"9C",x"5D",x"30",x"C9",x"19",x"80",x"A8",x"19", -- 0x3C88
		x"F5",x"06",x"BE",x"08",x"92",x"88",x"C9",x"2A", -- 0x3C90
		x"97",x"21",x"F1",x"3D",x"43",x"3E",x"7A",x"D0", -- 0x3C98
		x"E0",x"ED",x"AC",x"83",x"AE",x"D1",x"1F",x"0B", -- 0x3CA0
		x"62",x"20",x"96",x"78",x"B9",x"0B",x"49",x"08", -- 0x3CA8
		x"26",x"74",x"EE",x"F8",x"53",x"60",x"4D",x"17", -- 0x3CB0
		x"AD",x"85",x"59",x"54",x"E7",x"80",x"85",x"79", -- 0x3CB8
		x"1D",x"A5",x"29",x"A2",x"47",x"1A",x"84",x"11", -- 0x3CC0
		x"4C",x"A1",x"B6",x"80",x"FD",x"07",x"54",x"C5", -- 0x3CC8
		x"F1",x"46",x"5F",x"56",x"6A",x"36",x"56",x"93", -- 0x3CD0
		x"D3",x"29",x"7E",x"C4",x"37",x"CD",x"A5",x"49", -- 0x3CD8
		x"04",x"23",x"20",x"09",x"05",x"68",x"78",x"D9", -- 0x3CE0
		x"A7",x"C9",x"95",x"36",x"86",x"CC",x"A6",x"9E", -- 0x3CE8
		x"E1",x"3C",x"BF",x"42",x"D7",x"4A",x"D3",x"D4", -- 0x3CF0
		x"B6",x"81",x"BF",x"73",x"94",x"00",x"AF",x"EE", -- 0x3CF8
		x"C4",x"85",x"CC",x"11",x"EB",x"21",x"81",x"14", -- 0x3D00
		x"2A",x"54",x"06",x"5B",x"E0",x"F4",x"34",x"84", -- 0x3D08
		x"BA",x"4C",x"9B",x"1B",x"FB",x"01",x"8F",x"7E", -- 0x3D10
		x"E1",x"08",x"52",x"2A",x"A6",x"4A",x"A7",x"AA", -- 0x3D18
		x"84",x"82",x"2B",x"0E",x"6F",x"24",x"4B",x"8C", -- 0x3D20
		x"AD",x"09",x"94",x"0E",x"EF",x"47",x"2D",x"67", -- 0x3D28
		x"7C",x"34",x"FD",x"0E",x"74",x"0E",x"2A",x"75", -- 0x3D30
		x"86",x"C2",x"E7",x"A5",x"3B",x"6B",x"97",x"A6", -- 0x3D38
		x"75",x"80",x"D2",x"08",x"52",x"04",x"7E",x"1F", -- 0x3D40
		x"C8",x"42",x"84",x"15",x"CE",x"00",x"F8",x"00", -- 0x3D48
		x"72",x"A3",x"4A",x"D9",x"CD",x"A0",x"6A",x"8E", -- 0x3D50
		x"7F",x"C5",x"ED",x"07",x"7F",x"EF",x"5B",x"64", -- 0x3D58
		x"54",x"28",x"21",x"50",x"12",x"D3",x"B4",x"30", -- 0x3D60
		x"F7",x"0A",x"08",x"BC",x"ED",x"85",x"5F",x"0E", -- 0x3D68
		x"D2",x"BB",x"B3",x"BA",x"97",x"6D",x"F4",x"72", -- 0x3D70
		x"26",x"45",x"A3",x"86",x"93",x"72",x"7B",x"19", -- 0x3D78
		x"C5",x"41",x"29",x"10",x"7A",x"90",x"A3",x"B1", -- 0x3D80
		x"29",x"48",x"FA",x"B5",x"0C",x"07",x"27",x"98", -- 0x3D88
		x"EB",x"69",x"DA",x"10",x"DC",x"62",x"9C",x"3F", -- 0x3D90
		x"EF",x"42",x"6C",x"3A",x"FB",x"DB",x"29",x"7A", -- 0x3D98
		x"23",x"39",x"FD",x"A8",x"22",x"C5",x"F6",x"30", -- 0x3DA0
		x"D1",x"F5",x"F5",x"39",x"FD",x"FB",x"F6",x"0A", -- 0x3DA8
		x"E1",x"DB",x"D0",x"A4",x"36",x"4F",x"7D",x"B7", -- 0x3DB0
		x"FB",x"A4",x"70",x"8B",x"5C",x"CB",x"F7",x"52", -- 0x3DB8
		x"B0",x"52",x"82",x"83",x"05",x"10",x"CA",x"22", -- 0x3DC0
		x"26",x"01",x"19",x"01",x"C2",x"25",x"5E",x"C0", -- 0x3DC8
		x"29",x"45",x"B7",x"A3",x"CD",x"A2",x"BF",x"BD", -- 0x3DD0
		x"74",x"27",x"B6",x"F0",x"BD",x"4E",x"89",x"CB", -- 0x3DD8
		x"D6",x"0A",x"C6",x"4E",x"59",x"0C",x"4C",x"F9", -- 0x3DE0
		x"94",x"F2",x"16",x"A5",x"6B",x"C1",x"93",x"25", -- 0x3DE8
		x"67",x"AB",x"33",x"AF",x"3B",x"6B",x"C7",x"C5", -- 0x3DF0
		x"F5",x"1B",x"86",x"A8",x"F7",x"2C",x"CE",x"55", -- 0x3DF8
		x"37",x"01",x"47",x"07",x"45",x"16",x"12",x"00", -- 0x3E00
		x"49",x"89",x"B0",x"8A",x"48",x"02",x"63",x"CD", -- 0x3E08
		x"B3",x"01",x"99",x"59",x"B1",x"48",x"74",x"11", -- 0x3E10
		x"53",x"60",x"B0",x"2E",x"25",x"83",x"A5",x"74", -- 0x3E18
		x"7A",x"9D",x"0A",x"76",x"28",x"0D",x"7F",x"A4", -- 0x3E20
		x"B6",x"04",x"E6",x"AA",x"1F",x"25",x"9B",x"C4", -- 0x3E28
		x"F7",x"02",x"92",x"D2",x"44",x"EB",x"4B",x"0A", -- 0x3E30
		x"A3",x"8E",x"47",x"0E",x"D2",x"D0",x"8E",x"F9", -- 0x3E38
		x"AC",x"AD",x"01",x"08",x"3A",x"10",x"A7",x"22", -- 0x3E40
		x"30",x"C8",x"38",x"51",x"1B",x"C7",x"32",x"21", -- 0x3E48
		x"13",x"E2",x"4E",x"60",x"EC",x"E5",x"95",x"98", -- 0x3E50
		x"EC",x"02",x"4B",x"3D",x"65",x"A6",x"6A",x"D0", -- 0x3E58
		x"AD",x"77",x"97",x"51",x"82",x"68",x"4D",x"9B", -- 0x3E60
		x"9F",x"ED",x"7D",x"01",x"21",x"9F",x"EF",x"09", -- 0x3E68
		x"B8",x"7B",x"63",x"CA",x"FB",x"A3",x"87",x"4A", -- 0x3E70
		x"30",x"A5",x"86",x"FC",x"1F",x"E6",x"33",x"D7", -- 0x3E78
		x"FE",x"C1",x"96",x"59",x"8D",x"0B",x"BA",x"44", -- 0x3E80
		x"39",x"2A",x"73",x"0D",x"60",x"BC",x"D0",x"76", -- 0x3E88
		x"F5",x"55",x"BD",x"09",x"E5",x"91",x"48",x"52", -- 0x3E90
		x"22",x"00",x"9F",x"A3",x"8E",x"02",x"98",x"C1", -- 0x3E98
		x"0F",x"08",x"74",x"50",x"B7",x"AC",x"C6",x"80", -- 0x3EA0
		x"D4",x"81",x"6A",x"0F",x"D3",x"28",x"FD",x"49", -- 0x3EA8
		x"DC",x"04",x"5F",x"10",x"AF",x"87",x"76",x"06", -- 0x3EB0
		x"74",x"E6",x"E4",x"20",x"CB",x"A6",x"36",x"56", -- 0x3EB8
		x"3C",x"1E",x"4D",x"F2",x"03",x"06",x"9A",x"01", -- 0x3EC0
		x"C2",x"41",x"C9",x"01",x"D1",x"B5",x"10",x"30", -- 0x3EC8
		x"23",x"80",x"F2",x"0A",x"46",x"99",x"E7",x"22", -- 0x3ED0
		x"16",x"97",x"1A",x"48",x"10",x"A7",x"23",x"98", -- 0x3ED8
		x"DE",x"81",x"7C",x"23",x"F0",x"1F",x"14",x"33", -- 0x3EE0
		x"A3",x"94",x"CB",x"6D",x"59",x"CA",x"7B",x"9E", -- 0x3EE8
		x"1D",x"10",x"1F",x"C7",x"54",x"63",x"A4",x"0C", -- 0x3EF0
		x"F2",x"8C",x"93",x"0C",x"EA",x"78",x"AB",x"55", -- 0x3EF8
		x"C1",x"11",x"13",x"34",x"F1",x"05",x"74",x"22", -- 0x3F00
		x"BD",x"F0",x"6D",x"E5",x"38",x"10",x"16",x"30", -- 0x3F08
		x"1E",x"54",x"35",x"A6",x"9E",x"0D",x"E4",x"02", -- 0x3F10
		x"89",x"C5",x"8D",x"48",x"B0",x"34",x"F9",x"D0", -- 0x3F18
		x"54",x"07",x"7E",x"4A",x"91",x"06",x"88",x"22", -- 0x3F20
		x"43",x"3F",x"6B",x"50",x"6B",x"95",x"91",x"00", -- 0x3F28
		x"F9",x"A0",x"97",x"F5",x"8F",x"55",x"A5",x"49", -- 0x3F30
		x"3F",x"5B",x"51",x"6B",x"F4",x"38",x"F1",x"30", -- 0x3F38
		x"A2",x"00",x"45",x"81",x"49",x"4E",x"B8",x"58", -- 0x3F40
		x"49",x"A8",x"57",x"83",x"8B",x"E5",x"53",x"48", -- 0x3F48
		x"F9",x"9C",x"EE",x"90",x"5A",x"E5",x"D6",x"80", -- 0x3F50
		x"FF",x"74",x"B7",x"E1",x"FA",x"46",x"F1",x"15", -- 0x3F58
		x"B3",x"87",x"F2",x"BE",x"FD",x"21",x"7E",x"08", -- 0x3F60
		x"F7",x"D4",x"D7",x"E5",x"E7",x"40",x"12",x"C6", -- 0x3F68
		x"C1",x"9C",x"4D",x"0E",x"16",x"7D",x"32",x"09", -- 0x3F70
		x"57",x"10",x"BA",x"71",x"58",x"C7",x"F5",x"C0", -- 0x3F78
		x"EF",x"E4",x"FA",x"98",x"63",x"00",x"4D",x"8C", -- 0x3F80
		x"70",x"25",x"D2",x"12",x"DB",x"95",x"E3",x"C1", -- 0x3F88
		x"F0",x"1C",x"26",x"76",x"91",x"E0",x"47",x"AF", -- 0x3F90
		x"03",x"41",x"C9",x"06",x"24",x"98",x"72",x"2C", -- 0x3F98
		x"A6",x"8D",x"63",x"33",x"49",x"94",x"FD",x"B7", -- 0x3FA0
		x"C3",x"F8",x"65",x"A4",x"49",x"5A",x"2F",x"86", -- 0x3FA8
		x"8B",x"93",x"EB",x"43",x"1D",x"6A",x"6F",x"8C", -- 0x3FB0
		x"88",x"11",x"0A",x"88",x"AF",x"49",x"0D",x"42", -- 0x3FB8
		x"B9",x"72",x"30",x"0B",x"37",x"0F",x"83",x"18", -- 0x3FC0
		x"40",x"19",x"26",x"B7",x"B7",x"00",x"AB",x"92", -- 0x3FC8
		x"DB",x"F8",x"F5",x"00",x"DC",x"92",x"83",x"16", -- 0x3FD0
		x"83",x"B2",x"9B",x"53",x"F2",x"FC",x"4F",x"33", -- 0x3FD8
		x"79",x"CA",x"0C",x"C9",x"9F",x"E3",x"73",x"70", -- 0x3FE0
		x"67",x"A2",x"5C",x"A5",x"62",x"90",x"55",x"B7", -- 0x3FE8
		x"C9",x"81",x"6C",x"41",x"8F",x"67",x"3B",x"F6", -- 0x3FF0
		x"50",x"44",x"4E",x"3C",x"B1",x"38",x"47",x"42"  -- 0x3FF8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
  			DATA <= ROM(to_integer(unsigned(ADDR)));
		end if;
	end process;
end RTL;
